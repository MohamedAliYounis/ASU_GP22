module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;


 tile tile (.clk(wb_clk_i),
    .dyn0_dEo_valid(io_out[1]),
    .dyn0_dNo_valid(io_out[0]),
    .dyn0_dSo_valid(io_out[3]),
    .dyn0_dWo_valid(io_out[2]),
    .dyn0_yummyOut_E(io_out[5]),
    .dyn0_yummyOut_N(io_out[4]),
    .dyn0_yummyOut_S(io_out[7]),
    .dyn0_yummyOut_W(io_out[6]),
    .dyn1_dEo_valid(io_out[9]),
    .dyn1_dNo_valid(io_out[8]),
    .dyn1_dSo_valid(io_out[11]),
    .dyn1_dWo_valid(io_out[10]),
    .dyn1_yummyOut_E(io_out[13]),
    .dyn1_yummyOut_N(io_out[12]),
    .dyn1_yummyOut_S(io_out[15]),
    .dyn1_yummyOut_W(io_out[14]),
    .dyn2_dEo_valid(io_out[17]),
    .dyn2_dNo_valid(io_out[16]),
    .dyn2_dSo_valid(io_out[19]),
    .dyn2_dWo_valid(io_out[18]),
    .dyn2_yummyOut_E(io_out[21]),
    .dyn2_yummyOut_N(io_out[20]),
    .dyn2_yummyOut_S(io_out[23]),
    .dyn2_yummyOut_W(io_out[22]),
    .rst_n(wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .buffer_processor_data_noc1({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32,
    _NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40,
    _NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56,
    _NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .buffer_processor_data_noc3({_NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70,
    _NC71,
    _NC72,
    _NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80,
    _NC81,
    _NC82,
    _NC83,
    _NC84,
    _NC85,
    _NC86,
    _NC87,
    _NC88,
    _NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96,
    _NC97,
    _NC98,
    _NC99,
    _NC100,
    _NC101,
    _NC102,
    _NC103,
    _NC104,
    _NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112,
    _NC113,
    _NC114,
    _NC115,
    _NC116,
    _NC117,
    _NC118,
    _NC119,
    _NC120,
    _NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .chipid({_NC129,
    _NC130,
    _NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136,
    _NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142}),
    .config_chipid({_NC143,
    _NC144,
    _NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152,
    _NC153,
    _NC154,
    _NC155,
    _NC156}),
    .config_coreid_x({_NC157,
    _NC158,
    _NC159,
    _NC160,
    _NC161,
    _NC162,
    _NC163,
    _NC164}),
    .config_coreid_y({_NC165,
    _NC166,
    _NC167,
    _NC168,
    _NC169,
    _NC170,
    _NC171,
    _NC172}),
    .config_hmt_base({_NC173,
    _NC174,
    _NC175,
    _NC176,
    _NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184,
    _NC185,
    _NC186,
    _NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192,
    _NC193,
    _NC194}),
    .config_home_alloc_method({_NC195,
    _NC196}),
    .config_l15_read_res_data_s3({_NC197,
    _NC198,
    _NC199,
    _NC200,
    _NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208,
    _NC209,
    _NC210,
    _NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216,
    _NC217,
    _NC218,
    _NC219,
    _NC220,
    _NC221,
    _NC222,
    _NC223,
    _NC224,
    _NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232,
    _NC233,
    _NC234,
    _NC235,
    _NC236,
    _NC237,
    _NC238,
    _NC239,
    _NC240,
    _NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246,
    _NC247,
    _NC248,
    _NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256,
    _NC257,
    _NC258,
    _NC259,
    _NC260}),
    .config_system_tile_count_5_0({_NC261,
    _NC262,
    _NC263,
    _NC264,
    _NC265,
    _NC266}),
    .coreid_x({_NC267,
    _NC268,
    _NC269,
    _NC270,
    _NC271,
    _NC272,
    _NC273,
    _NC274}),
    .coreid_y({_NC275,
    _NC276,
    _NC277,
    _NC278,
    _NC279,
    _NC280,
    _NC281,
    _NC282}),
    .default_chipid({_NC283,
    _NC284,
    _NC285,
    _NC286,
    _NC287,
    _NC288,
    _NC289,
    _NC290,
    _NC291,
    _NC292,
    _NC293,
    _NC294,
    _NC295,
    _NC296}),
    .default_coreid_x({_NC297,
    _NC298,
    _NC299,
    _NC300,
    _NC301,
    _NC302,
    _NC303,
    _NC304}),
    .default_coreid_y({_NC305,
    _NC306,
    _NC307,
    _NC308,
    _NC309,
    _NC310,
    _NC311,
    _NC312}),
    .dummy_core({_NC313,
    _NC314,
    _NC315,
    _NC316,
    _NC317,
    _NC318,
    _NC319,
    _NC320,
    _NC321,
    _NC322,
    _NC323,
    _NC324,
    _NC325,
    _NC326,
    _NC327,
    _NC328,
    _NC329,
    _NC330,
    _NC331,
    _NC332,
    _NC333,
    _NC334,
    _NC335,
    _NC336,
    _NC337,
    _NC338,
    _NC339,
    _NC340,
    _NC341,
    _NC342,
    _NC343,
    _NC344}),
    .dyn0_dEo({_NC345,
    _NC346,
    _NC347,
    _NC348,
    _NC349,
    _NC350,
    _NC351,
    _NC352,
    _NC353,
    _NC354,
    _NC355,
    _NC356,
    _NC357,
    _NC358,
    _NC359,
    _NC360,
    _NC361,
    _NC362,
    _NC363,
    _NC364,
    _NC365,
    _NC366,
    _NC367,
    _NC368,
    _NC369,
    _NC370,
    _NC371,
    _NC372,
    _NC373,
    _NC374,
    _NC375,
    _NC376,
    _NC377,
    _NC378,
    _NC379,
    _NC380,
    _NC381,
    _NC382,
    _NC383,
    _NC384,
    _NC385,
    _NC386,
    _NC387,
    _NC388,
    _NC389,
    _NC390,
    _NC391,
    _NC392,
    _NC393,
    _NC394,
    _NC395,
    _NC396,
    _NC397,
    _NC398,
    _NC399,
    _NC400,
    _NC401,
    _NC402,
    _NC403,
    _NC404,
    _NC405,
    _NC406,
    _NC407,
    _NC408}),
    .dyn0_dNo({_NC409,
    _NC410,
    _NC411,
    _NC412,
    _NC413,
    _NC414,
    _NC415,
    _NC416,
    _NC417,
    _NC418,
    _NC419,
    _NC420,
    _NC421,
    _NC422,
    _NC423,
    _NC424,
    _NC425,
    _NC426,
    _NC427,
    _NC428,
    _NC429,
    _NC430,
    _NC431,
    _NC432,
    _NC433,
    _NC434,
    _NC435,
    _NC436,
    _NC437,
    _NC438,
    _NC439,
    _NC440,
    _NC441,
    _NC442,
    _NC443,
    _NC444,
    _NC445,
    _NC446,
    _NC447,
    _NC448,
    _NC449,
    _NC450,
    _NC451,
    _NC452,
    _NC453,
    _NC454,
    _NC455,
    _NC456,
    _NC457,
    _NC458,
    _NC459,
    _NC460,
    _NC461,
    _NC462,
    _NC463,
    _NC464,
    _NC465,
    _NC466,
    _NC467,
    _NC468,
    _NC469,
    _NC470,
    _NC471,
    _NC472}),
    .dyn0_dSo({_NC473,
    _NC474,
    _NC475,
    _NC476,
    _NC477,
    _NC478,
    _NC479,
    _NC480,
    _NC481,
    _NC482,
    _NC483,
    _NC484,
    _NC485,
    _NC486,
    _NC487,
    _NC488,
    _NC489,
    _NC490,
    _NC491,
    _NC492,
    _NC493,
    _NC494,
    _NC495,
    _NC496,
    _NC497,
    _NC498,
    _NC499,
    _NC500,
    _NC501,
    _NC502,
    _NC503,
    _NC504,
    _NC505,
    _NC506,
    _NC507,
    _NC508,
    _NC509,
    _NC510,
    _NC511,
    _NC512,
    _NC513,
    _NC514,
    _NC515,
    _NC516,
    _NC517,
    _NC518,
    _NC519,
    _NC520,
    _NC521,
    _NC522,
    _NC523,
    _NC524,
    _NC525,
    _NC526,
    _NC527,
    _NC528,
    _NC529,
    _NC530,
    _NC531,
    _NC532,
    _NC533,
    _NC534,
    _NC535,
    _NC536}),
    .dyn0_dWo({_NC537,
    _NC538,
    _NC539,
    _NC540,
    _NC541,
    _NC542,
    _NC543,
    _NC544,
    _NC545,
    _NC546,
    _NC547,
    _NC548,
    _NC549,
    _NC550,
    _NC551,
    _NC552,
    _NC553,
    _NC554,
    _NC555,
    _NC556,
    _NC557,
    _NC558,
    _NC559,
    _NC560,
    _NC561,
    _NC562,
    _NC563,
    _NC564,
    _NC565,
    _NC566,
    _NC567,
    _NC568,
    _NC569,
    _NC570,
    _NC571,
    _NC572,
    _NC573,
    _NC574,
    _NC575,
    _NC576,
    _NC577,
    _NC578,
    _NC579,
    _NC580,
    _NC581,
    _NC582,
    _NC583,
    _NC584,
    _NC585,
    _NC586,
    _NC587,
    _NC588,
    _NC589,
    _NC590,
    _NC591,
    _NC592,
    _NC593,
    _NC594,
    _NC595,
    _NC596,
    _NC597,
    _NC598,
    _NC599,
    _NC600}),
    .dyn0_dataIn_E({_NC601,
    _NC602,
    _NC603,
    _NC604,
    _NC605,
    _NC606,
    _NC607,
    _NC608,
    _NC609,
    _NC610,
    _NC611,
    _NC612,
    _NC613,
    _NC614,
    _NC615,
    _NC616,
    _NC617,
    _NC618,
    _NC619,
    _NC620,
    _NC621,
    _NC622,
    _NC623,
    _NC624,
    _NC625,
    _NC626,
    _NC627,
    _NC628,
    _NC629,
    _NC630,
    _NC631,
    _NC632,
    _NC633,
    _NC634,
    _NC635,
    _NC636,
    _NC637,
    _NC638,
    _NC639,
    _NC640,
    _NC641,
    _NC642,
    _NC643,
    _NC644,
    _NC645,
    _NC646,
    _NC647,
    _NC648,
    _NC649,
    _NC650,
    _NC651,
    _NC652,
    _NC653,
    _NC654,
    _NC655,
    _NC656,
    _NC657,
    _NC658,
    _NC659,
    _NC660,
    _NC661,
    _NC662,
    _NC663,
    _NC664}),
    .dyn0_dataIn_N({_NC665,
    _NC666,
    _NC667,
    _NC668,
    _NC669,
    _NC670,
    _NC671,
    _NC672,
    _NC673,
    _NC674,
    _NC675,
    _NC676,
    _NC677,
    _NC678,
    _NC679,
    _NC680,
    _NC681,
    _NC682,
    _NC683,
    _NC684,
    _NC685,
    _NC686,
    _NC687,
    _NC688,
    _NC689,
    _NC690,
    _NC691,
    _NC692,
    _NC693,
    _NC694,
    _NC695,
    _NC696,
    _NC697,
    _NC698,
    _NC699,
    _NC700,
    _NC701,
    _NC702,
    _NC703,
    _NC704,
    _NC705,
    _NC706,
    _NC707,
    _NC708,
    _NC709,
    _NC710,
    _NC711,
    _NC712,
    _NC713,
    _NC714,
    _NC715,
    _NC716,
    _NC717,
    _NC718,
    _NC719,
    _NC720,
    _NC721,
    _NC722,
    _NC723,
    _NC724,
    _NC725,
    _NC726,
    _NC727,
    _NC728}),
    .dyn0_dataIn_S({_NC729,
    _NC730,
    _NC731,
    _NC732,
    _NC733,
    _NC734,
    _NC735,
    _NC736,
    _NC737,
    _NC738,
    _NC739,
    _NC740,
    _NC741,
    _NC742,
    _NC743,
    _NC744,
    _NC745,
    _NC746,
    _NC747,
    _NC748,
    _NC749,
    _NC750,
    _NC751,
    _NC752,
    _NC753,
    _NC754,
    _NC755,
    _NC756,
    _NC757,
    _NC758,
    _NC759,
    _NC760,
    _NC761,
    _NC762,
    _NC763,
    _NC764,
    _NC765,
    _NC766,
    _NC767,
    _NC768,
    _NC769,
    _NC770,
    _NC771,
    _NC772,
    _NC773,
    _NC774,
    _NC775,
    _NC776,
    _NC777,
    _NC778,
    _NC779,
    _NC780,
    _NC781,
    _NC782,
    _NC783,
    _NC784,
    _NC785,
    _NC786,
    _NC787,
    _NC788,
    _NC789,
    _NC790,
    _NC791,
    _NC792}),
    .dyn0_dataIn_W({_NC793,
    _NC794,
    _NC795,
    _NC796,
    _NC797,
    _NC798,
    _NC799,
    _NC800,
    _NC801,
    _NC802,
    _NC803,
    _NC804,
    _NC805,
    _NC806,
    _NC807,
    _NC808,
    _NC809,
    _NC810,
    _NC811,
    _NC812,
    _NC813,
    _NC814,
    _NC815,
    _NC816,
    _NC817,
    _NC818,
    _NC819,
    _NC820,
    _NC821,
    _NC822,
    _NC823,
    _NC824,
    _NC825,
    _NC826,
    _NC827,
    _NC828,
    _NC829,
    _NC830,
    _NC831,
    _NC832,
    _NC833,
    _NC834,
    _NC835,
    _NC836,
    _NC837,
    _NC838,
    _NC839,
    _NC840,
    _NC841,
    _NC842,
    _NC843,
    _NC844,
    _NC845,
    _NC846,
    _NC847,
    _NC848,
    _NC849,
    _NC850,
    _NC851,
    _NC852,
    _NC853,
    _NC854,
    _NC855,
    _NC856}),
    .dyn1_dEo({_NC857,
    _NC858,
    _NC859,
    _NC860,
    _NC861,
    _NC862,
    _NC863,
    _NC864,
    _NC865,
    _NC866,
    _NC867,
    _NC868,
    _NC869,
    _NC870,
    _NC871,
    _NC872,
    _NC873,
    _NC874,
    _NC875,
    _NC876,
    _NC877,
    _NC878,
    _NC879,
    _NC880,
    _NC881,
    _NC882,
    _NC883,
    _NC884,
    _NC885,
    _NC886,
    _NC887,
    _NC888,
    _NC889,
    _NC890,
    _NC891,
    _NC892,
    _NC893,
    _NC894,
    _NC895,
    _NC896,
    _NC897,
    _NC898,
    _NC899,
    _NC900,
    _NC901,
    _NC902,
    _NC903,
    _NC904,
    _NC905,
    _NC906,
    _NC907,
    _NC908,
    _NC909,
    _NC910,
    _NC911,
    _NC912,
    _NC913,
    _NC914,
    _NC915,
    _NC916,
    _NC917,
    _NC918,
    _NC919,
    _NC920}),
    .dyn1_dNo({_NC921,
    _NC922,
    _NC923,
    _NC924,
    _NC925,
    _NC926,
    _NC927,
    _NC928,
    _NC929,
    _NC930,
    _NC931,
    _NC932,
    _NC933,
    _NC934,
    _NC935,
    _NC936,
    _NC937,
    _NC938,
    _NC939,
    _NC940,
    _NC941,
    _NC942,
    _NC943,
    _NC944,
    _NC945,
    _NC946,
    _NC947,
    _NC948,
    _NC949,
    _NC950,
    _NC951,
    _NC952,
    _NC953,
    _NC954,
    _NC955,
    _NC956,
    _NC957,
    _NC958,
    _NC959,
    _NC960,
    _NC961,
    _NC962,
    _NC963,
    _NC964,
    _NC965,
    _NC966,
    _NC967,
    _NC968,
    _NC969,
    _NC970,
    _NC971,
    _NC972,
    _NC973,
    _NC974,
    _NC975,
    _NC976,
    _NC977,
    _NC978,
    _NC979,
    _NC980,
    _NC981,
    _NC982,
    _NC983,
    _NC984}),
    .dyn1_dSo({_NC985,
    _NC986,
    _NC987,
    _NC988,
    _NC989,
    _NC990,
    _NC991,
    _NC992,
    _NC993,
    _NC994,
    _NC995,
    _NC996,
    _NC997,
    _NC998,
    _NC999,
    _NC1000,
    _NC1001,
    _NC1002,
    _NC1003,
    _NC1004,
    _NC1005,
    _NC1006,
    _NC1007,
    _NC1008,
    _NC1009,
    _NC1010,
    _NC1011,
    _NC1012,
    _NC1013,
    _NC1014,
    _NC1015,
    _NC1016,
    _NC1017,
    _NC1018,
    _NC1019,
    _NC1020,
    _NC1021,
    _NC1022,
    _NC1023,
    _NC1024,
    _NC1025,
    _NC1026,
    _NC1027,
    _NC1028,
    _NC1029,
    _NC1030,
    _NC1031,
    _NC1032,
    _NC1033,
    _NC1034,
    _NC1035,
    _NC1036,
    _NC1037,
    _NC1038,
    _NC1039,
    _NC1040,
    _NC1041,
    _NC1042,
    _NC1043,
    _NC1044,
    _NC1045,
    _NC1046,
    _NC1047,
    _NC1048}),
    .dyn1_dWo({_NC1049,
    _NC1050,
    _NC1051,
    _NC1052,
    _NC1053,
    _NC1054,
    _NC1055,
    _NC1056,
    _NC1057,
    _NC1058,
    _NC1059,
    _NC1060,
    _NC1061,
    _NC1062,
    _NC1063,
    _NC1064,
    _NC1065,
    _NC1066,
    _NC1067,
    _NC1068,
    _NC1069,
    _NC1070,
    _NC1071,
    _NC1072,
    _NC1073,
    _NC1074,
    _NC1075,
    _NC1076,
    _NC1077,
    _NC1078,
    _NC1079,
    _NC1080,
    _NC1081,
    _NC1082,
    _NC1083,
    _NC1084,
    _NC1085,
    _NC1086,
    _NC1087,
    _NC1088,
    _NC1089,
    _NC1090,
    _NC1091,
    _NC1092,
    _NC1093,
    _NC1094,
    _NC1095,
    _NC1096,
    _NC1097,
    _NC1098,
    _NC1099,
    _NC1100,
    _NC1101,
    _NC1102,
    _NC1103,
    _NC1104,
    _NC1105,
    _NC1106,
    _NC1107,
    _NC1108,
    _NC1109,
    _NC1110,
    _NC1111,
    _NC1112}),
    .dyn1_dataIn_E({_NC1113,
    _NC1114,
    _NC1115,
    _NC1116,
    _NC1117,
    _NC1118,
    _NC1119,
    _NC1120,
    _NC1121,
    _NC1122,
    _NC1123,
    _NC1124,
    _NC1125,
    _NC1126,
    _NC1127,
    _NC1128,
    _NC1129,
    _NC1130,
    _NC1131,
    _NC1132,
    _NC1133,
    _NC1134,
    _NC1135,
    _NC1136,
    _NC1137,
    _NC1138,
    _NC1139,
    _NC1140,
    _NC1141,
    _NC1142,
    _NC1143,
    _NC1144,
    _NC1145,
    _NC1146,
    _NC1147,
    _NC1148,
    _NC1149,
    _NC1150,
    _NC1151,
    _NC1152,
    _NC1153,
    _NC1154,
    _NC1155,
    _NC1156,
    _NC1157,
    _NC1158,
    _NC1159,
    _NC1160,
    _NC1161,
    _NC1162,
    _NC1163,
    _NC1164,
    _NC1165,
    _NC1166,
    _NC1167,
    _NC1168,
    _NC1169,
    _NC1170,
    _NC1171,
    _NC1172,
    _NC1173,
    _NC1174,
    _NC1175,
    _NC1176}),
    .dyn1_dataIn_N({_NC1177,
    _NC1178,
    _NC1179,
    _NC1180,
    _NC1181,
    _NC1182,
    _NC1183,
    _NC1184,
    _NC1185,
    _NC1186,
    _NC1187,
    _NC1188,
    _NC1189,
    _NC1190,
    _NC1191,
    _NC1192,
    _NC1193,
    _NC1194,
    _NC1195,
    _NC1196,
    _NC1197,
    _NC1198,
    _NC1199,
    _NC1200,
    _NC1201,
    _NC1202,
    _NC1203,
    _NC1204,
    _NC1205,
    _NC1206,
    _NC1207,
    _NC1208,
    _NC1209,
    _NC1210,
    _NC1211,
    _NC1212,
    _NC1213,
    _NC1214,
    _NC1215,
    _NC1216,
    _NC1217,
    _NC1218,
    _NC1219,
    _NC1220,
    _NC1221,
    _NC1222,
    _NC1223,
    _NC1224,
    _NC1225,
    _NC1226,
    _NC1227,
    _NC1228,
    _NC1229,
    _NC1230,
    _NC1231,
    _NC1232,
    _NC1233,
    _NC1234,
    _NC1235,
    _NC1236,
    _NC1237,
    _NC1238,
    _NC1239,
    _NC1240}),
    .dyn1_dataIn_S({_NC1241,
    _NC1242,
    _NC1243,
    _NC1244,
    _NC1245,
    _NC1246,
    _NC1247,
    _NC1248,
    _NC1249,
    _NC1250,
    _NC1251,
    _NC1252,
    _NC1253,
    _NC1254,
    _NC1255,
    _NC1256,
    _NC1257,
    _NC1258,
    _NC1259,
    _NC1260,
    _NC1261,
    _NC1262,
    _NC1263,
    _NC1264,
    _NC1265,
    _NC1266,
    _NC1267,
    _NC1268,
    _NC1269,
    _NC1270,
    _NC1271,
    _NC1272,
    _NC1273,
    _NC1274,
    _NC1275,
    _NC1276,
    _NC1277,
    _NC1278,
    _NC1279,
    _NC1280,
    _NC1281,
    _NC1282,
    _NC1283,
    _NC1284,
    _NC1285,
    _NC1286,
    _NC1287,
    _NC1288,
    _NC1289,
    _NC1290,
    _NC1291,
    _NC1292,
    _NC1293,
    _NC1294,
    _NC1295,
    _NC1296,
    _NC1297,
    _NC1298,
    _NC1299,
    _NC1300,
    _NC1301,
    _NC1302,
    _NC1303,
    _NC1304}),
    .dyn1_dataIn_W({_NC1305,
    _NC1306,
    _NC1307,
    _NC1308,
    _NC1309,
    _NC1310,
    _NC1311,
    _NC1312,
    _NC1313,
    _NC1314,
    _NC1315,
    _NC1316,
    _NC1317,
    _NC1318,
    _NC1319,
    _NC1320,
    _NC1321,
    _NC1322,
    _NC1323,
    _NC1324,
    _NC1325,
    _NC1326,
    _NC1327,
    _NC1328,
    _NC1329,
    _NC1330,
    _NC1331,
    _NC1332,
    _NC1333,
    _NC1334,
    _NC1335,
    _NC1336,
    _NC1337,
    _NC1338,
    _NC1339,
    _NC1340,
    _NC1341,
    _NC1342,
    _NC1343,
    _NC1344,
    _NC1345,
    _NC1346,
    _NC1347,
    _NC1348,
    _NC1349,
    _NC1350,
    _NC1351,
    _NC1352,
    _NC1353,
    _NC1354,
    _NC1355,
    _NC1356,
    _NC1357,
    _NC1358,
    _NC1359,
    _NC1360,
    _NC1361,
    _NC1362,
    _NC1363,
    _NC1364,
    _NC1365,
    _NC1366,
    _NC1367,
    _NC1368}),
    .dyn2_dEo({_NC1369,
    _NC1370,
    _NC1371,
    _NC1372,
    _NC1373,
    _NC1374,
    _NC1375,
    _NC1376,
    _NC1377,
    _NC1378,
    _NC1379,
    _NC1380,
    _NC1381,
    _NC1382,
    _NC1383,
    _NC1384,
    _NC1385,
    _NC1386,
    _NC1387,
    _NC1388,
    _NC1389,
    _NC1390,
    _NC1391,
    _NC1392,
    _NC1393,
    _NC1394,
    _NC1395,
    _NC1396,
    _NC1397,
    _NC1398,
    _NC1399,
    _NC1400,
    _NC1401,
    _NC1402,
    _NC1403,
    _NC1404,
    _NC1405,
    _NC1406,
    _NC1407,
    _NC1408,
    _NC1409,
    _NC1410,
    _NC1411,
    _NC1412,
    _NC1413,
    _NC1414,
    _NC1415,
    _NC1416,
    _NC1417,
    _NC1418,
    _NC1419,
    _NC1420,
    _NC1421,
    _NC1422,
    _NC1423,
    _NC1424,
    _NC1425,
    _NC1426,
    _NC1427,
    _NC1428,
    _NC1429,
    _NC1430,
    _NC1431,
    _NC1432}),
    .dyn2_dNo({_NC1433,
    _NC1434,
    _NC1435,
    _NC1436,
    _NC1437,
    _NC1438,
    _NC1439,
    _NC1440,
    _NC1441,
    _NC1442,
    _NC1443,
    _NC1444,
    _NC1445,
    _NC1446,
    _NC1447,
    _NC1448,
    _NC1449,
    _NC1450,
    _NC1451,
    _NC1452,
    _NC1453,
    _NC1454,
    _NC1455,
    _NC1456,
    _NC1457,
    _NC1458,
    _NC1459,
    _NC1460,
    _NC1461,
    _NC1462,
    _NC1463,
    _NC1464,
    _NC1465,
    _NC1466,
    _NC1467,
    _NC1468,
    _NC1469,
    _NC1470,
    _NC1471,
    _NC1472,
    _NC1473,
    _NC1474,
    _NC1475,
    _NC1476,
    _NC1477,
    _NC1478,
    _NC1479,
    _NC1480,
    _NC1481,
    _NC1482,
    _NC1483,
    _NC1484,
    _NC1485,
    _NC1486,
    _NC1487,
    _NC1488,
    _NC1489,
    _NC1490,
    _NC1491,
    _NC1492,
    _NC1493,
    _NC1494,
    _NC1495,
    _NC1496}),
    .dyn2_dSo({_NC1497,
    _NC1498,
    _NC1499,
    _NC1500,
    _NC1501,
    _NC1502,
    _NC1503,
    _NC1504,
    _NC1505,
    _NC1506,
    _NC1507,
    _NC1508,
    _NC1509,
    _NC1510,
    _NC1511,
    _NC1512,
    _NC1513,
    _NC1514,
    _NC1515,
    _NC1516,
    _NC1517,
    _NC1518,
    _NC1519,
    _NC1520,
    _NC1521,
    _NC1522,
    _NC1523,
    _NC1524,
    _NC1525,
    _NC1526,
    _NC1527,
    _NC1528,
    _NC1529,
    _NC1530,
    _NC1531,
    _NC1532,
    _NC1533,
    _NC1534,
    _NC1535,
    _NC1536,
    _NC1537,
    _NC1538,
    _NC1539,
    _NC1540,
    _NC1541,
    _NC1542,
    _NC1543,
    _NC1544,
    _NC1545,
    _NC1546,
    _NC1547,
    _NC1548,
    _NC1549,
    _NC1550,
    _NC1551,
    _NC1552,
    _NC1553,
    _NC1554,
    _NC1555,
    _NC1556,
    _NC1557,
    _NC1558,
    _NC1559,
    _NC1560}),
    .dyn2_dWo({_NC1561,
    _NC1562,
    _NC1563,
    _NC1564,
    _NC1565,
    _NC1566,
    _NC1567,
    _NC1568,
    _NC1569,
    _NC1570,
    _NC1571,
    _NC1572,
    _NC1573,
    _NC1574,
    _NC1575,
    _NC1576,
    _NC1577,
    _NC1578,
    _NC1579,
    _NC1580,
    _NC1581,
    _NC1582,
    _NC1583,
    _NC1584,
    _NC1585,
    _NC1586,
    _NC1587,
    _NC1588,
    _NC1589,
    _NC1590,
    _NC1591,
    _NC1592,
    _NC1593,
    _NC1594,
    _NC1595,
    _NC1596,
    _NC1597,
    _NC1598,
    _NC1599,
    _NC1600,
    _NC1601,
    _NC1602,
    _NC1603,
    _NC1604,
    _NC1605,
    _NC1606,
    _NC1607,
    _NC1608,
    _NC1609,
    _NC1610,
    _NC1611,
    _NC1612,
    _NC1613,
    _NC1614,
    _NC1615,
    _NC1616,
    _NC1617,
    _NC1618,
    _NC1619,
    _NC1620,
    _NC1621,
    _NC1622,
    _NC1623,
    _NC1624}),
    .dyn2_dataIn_E({_NC1625,
    _NC1626,
    _NC1627,
    _NC1628,
    _NC1629,
    _NC1630,
    _NC1631,
    _NC1632,
    _NC1633,
    _NC1634,
    _NC1635,
    _NC1636,
    _NC1637,
    _NC1638,
    _NC1639,
    _NC1640,
    _NC1641,
    _NC1642,
    _NC1643,
    _NC1644,
    _NC1645,
    _NC1646,
    _NC1647,
    _NC1648,
    _NC1649,
    _NC1650,
    _NC1651,
    _NC1652,
    _NC1653,
    _NC1654,
    _NC1655,
    _NC1656,
    _NC1657,
    _NC1658,
    _NC1659,
    _NC1660,
    _NC1661,
    _NC1662,
    _NC1663,
    _NC1664,
    _NC1665,
    _NC1666,
    _NC1667,
    _NC1668,
    _NC1669,
    _NC1670,
    _NC1671,
    _NC1672,
    _NC1673,
    _NC1674,
    _NC1675,
    _NC1676,
    _NC1677,
    _NC1678,
    _NC1679,
    _NC1680,
    _NC1681,
    _NC1682,
    _NC1683,
    _NC1684,
    _NC1685,
    _NC1686,
    _NC1687,
    _NC1688}),
    .dyn2_dataIn_N({_NC1689,
    _NC1690,
    _NC1691,
    _NC1692,
    _NC1693,
    _NC1694,
    _NC1695,
    _NC1696,
    _NC1697,
    _NC1698,
    _NC1699,
    _NC1700,
    _NC1701,
    _NC1702,
    _NC1703,
    _NC1704,
    _NC1705,
    _NC1706,
    _NC1707,
    _NC1708,
    _NC1709,
    _NC1710,
    _NC1711,
    _NC1712,
    _NC1713,
    _NC1714,
    _NC1715,
    _NC1716,
    _NC1717,
    _NC1718,
    _NC1719,
    _NC1720,
    _NC1721,
    _NC1722,
    _NC1723,
    _NC1724,
    _NC1725,
    _NC1726,
    _NC1727,
    _NC1728,
    _NC1729,
    _NC1730,
    _NC1731,
    _NC1732,
    _NC1733,
    _NC1734,
    _NC1735,
    _NC1736,
    _NC1737,
    _NC1738,
    _NC1739,
    _NC1740,
    _NC1741,
    _NC1742,
    _NC1743,
    _NC1744,
    _NC1745,
    _NC1746,
    _NC1747,
    _NC1748,
    _NC1749,
    _NC1750,
    _NC1751,
    _NC1752}),
    .dyn2_dataIn_S({_NC1753,
    _NC1754,
    _NC1755,
    _NC1756,
    _NC1757,
    _NC1758,
    _NC1759,
    _NC1760,
    _NC1761,
    _NC1762,
    _NC1763,
    _NC1764,
    _NC1765,
    _NC1766,
    _NC1767,
    _NC1768,
    _NC1769,
    _NC1770,
    _NC1771,
    _NC1772,
    _NC1773,
    _NC1774,
    _NC1775,
    _NC1776,
    _NC1777,
    _NC1778,
    _NC1779,
    _NC1780,
    _NC1781,
    _NC1782,
    _NC1783,
    _NC1784,
    _NC1785,
    _NC1786,
    _NC1787,
    _NC1788,
    _NC1789,
    _NC1790,
    _NC1791,
    _NC1792,
    _NC1793,
    _NC1794,
    _NC1795,
    _NC1796,
    _NC1797,
    _NC1798,
    _NC1799,
    _NC1800,
    _NC1801,
    _NC1802,
    _NC1803,
    _NC1804,
    _NC1805,
    _NC1806,
    _NC1807,
    _NC1808,
    _NC1809,
    _NC1810,
    _NC1811,
    _NC1812,
    _NC1813,
    _NC1814,
    _NC1815,
    _NC1816}),
    .dyn2_dataIn_W({_NC1817,
    _NC1818,
    _NC1819,
    _NC1820,
    _NC1821,
    _NC1822,
    _NC1823,
    _NC1824,
    _NC1825,
    _NC1826,
    _NC1827,
    _NC1828,
    _NC1829,
    _NC1830,
    _NC1831,
    _NC1832,
    _NC1833,
    _NC1834,
    _NC1835,
    _NC1836,
    _NC1837,
    _NC1838,
    _NC1839,
    _NC1840,
    _NC1841,
    _NC1842,
    _NC1843,
    _NC1844,
    _NC1845,
    _NC1846,
    _NC1847,
    _NC1848,
    _NC1849,
    _NC1850,
    _NC1851,
    _NC1852,
    _NC1853,
    _NC1854,
    _NC1855,
    _NC1856,
    _NC1857,
    _NC1858,
    _NC1859,
    _NC1860,
    _NC1861,
    _NC1862,
    _NC1863,
    _NC1864,
    _NC1865,
    _NC1866,
    _NC1867,
    _NC1868,
    _NC1869,
    _NC1870,
    _NC1871,
    _NC1872,
    _NC1873,
    _NC1874,
    _NC1875,
    _NC1876,
    _NC1877,
    _NC1878,
    _NC1879,
    _NC1880}),
    .flat_tileid({_NC1881,
    _NC1882,
    _NC1883,
    _NC1884,
    _NC1885,
    _NC1886,
    _NC1887,
    _NC1888}),
    .jtag_tiles_ucb_data({_NC1889,
    _NC1890,
    _NC1891,
    _NC1892}),
    .l15_config_req_address_s2({_NC1893,
    _NC1894,
    _NC1895,
    _NC1896,
    _NC1897,
    _NC1898,
    _NC1899,
    _NC1900}),
    .l15_config_write_req_data_s2({_NC1901,
    _NC1902,
    _NC1903,
    _NC1904,
    _NC1905,
    _NC1906,
    _NC1907,
    _NC1908,
    _NC1909,
    _NC1910,
    _NC1911,
    _NC1912,
    _NC1913,
    _NC1914,
    _NC1915,
    _NC1916,
    _NC1917,
    _NC1918,
    _NC1919,
    _NC1920,
    _NC1921,
    _NC1922,
    _NC1923,
    _NC1924,
    _NC1925,
    _NC1926,
    _NC1927,
    _NC1928,
    _NC1929,
    _NC1930,
    _NC1931,
    _NC1932,
    _NC1933,
    _NC1934,
    _NC1935,
    _NC1936,
    _NC1937,
    _NC1938,
    _NC1939,
    _NC1940,
    _NC1941,
    _NC1942,
    _NC1943,
    _NC1944,
    _NC1945,
    _NC1946,
    _NC1947,
    _NC1948,
    _NC1949,
    _NC1950,
    _NC1951,
    _NC1952,
    _NC1953,
    _NC1954,
    _NC1955,
    _NC1956,
    _NC1957,
    _NC1958,
    _NC1959,
    _NC1960,
    _NC1961,
    _NC1962,
    _NC1963,
    _NC1964}),
    .l15_dmbr_l1missTag({_NC1965,
    _NC1966,
    _NC1967,
    _NC1968}),
    .l15_dmbr_l2missTag({_NC1969,
    _NC1970,
    _NC1971,
    _NC1972}),
    .l15_transducer_cross_invalidate_way({_NC1973,
    _NC1974}),
    .l15_transducer_data_0({_NC1975,
    _NC1976,
    _NC1977,
    _NC1978,
    _NC1979,
    _NC1980,
    _NC1981,
    _NC1982,
    _NC1983,
    _NC1984,
    _NC1985,
    _NC1986,
    _NC1987,
    _NC1988,
    _NC1989,
    _NC1990,
    _NC1991,
    _NC1992,
    _NC1993,
    _NC1994,
    _NC1995,
    _NC1996,
    _NC1997,
    _NC1998,
    _NC1999,
    _NC2000,
    _NC2001,
    _NC2002,
    _NC2003,
    _NC2004,
    _NC2005,
    _NC2006,
    _NC2007,
    _NC2008,
    _NC2009,
    _NC2010,
    _NC2011,
    _NC2012,
    _NC2013,
    _NC2014,
    _NC2015,
    _NC2016,
    _NC2017,
    _NC2018,
    _NC2019,
    _NC2020,
    _NC2021,
    _NC2022,
    _NC2023,
    _NC2024,
    _NC2025,
    _NC2026,
    _NC2027,
    _NC2028,
    _NC2029,
    _NC2030,
    _NC2031,
    _NC2032,
    _NC2033,
    _NC2034,
    _NC2035,
    _NC2036,
    _NC2037,
    _NC2038}),
    .l15_transducer_data_1({_NC2039,
    _NC2040,
    _NC2041,
    _NC2042,
    _NC2043,
    _NC2044,
    _NC2045,
    _NC2046,
    _NC2047,
    _NC2048,
    _NC2049,
    _NC2050,
    _NC2051,
    _NC2052,
    _NC2053,
    _NC2054,
    _NC2055,
    _NC2056,
    _NC2057,
    _NC2058,
    _NC2059,
    _NC2060,
    _NC2061,
    _NC2062,
    _NC2063,
    _NC2064,
    _NC2065,
    _NC2066,
    _NC2067,
    _NC2068,
    _NC2069,
    _NC2070,
    _NC2071,
    _NC2072,
    _NC2073,
    _NC2074,
    _NC2075,
    _NC2076,
    _NC2077,
    _NC2078,
    _NC2079,
    _NC2080,
    _NC2081,
    _NC2082,
    _NC2083,
    _NC2084,
    _NC2085,
    _NC2086,
    _NC2087,
    _NC2088,
    _NC2089,
    _NC2090,
    _NC2091,
    _NC2092,
    _NC2093,
    _NC2094,
    _NC2095,
    _NC2096,
    _NC2097,
    _NC2098,
    _NC2099,
    _NC2100,
    _NC2101,
    _NC2102}),
    .l15_transducer_data_2({_NC2103,
    _NC2104,
    _NC2105,
    _NC2106,
    _NC2107,
    _NC2108,
    _NC2109,
    _NC2110,
    _NC2111,
    _NC2112,
    _NC2113,
    _NC2114,
    _NC2115,
    _NC2116,
    _NC2117,
    _NC2118,
    _NC2119,
    _NC2120,
    _NC2121,
    _NC2122,
    _NC2123,
    _NC2124,
    _NC2125,
    _NC2126,
    _NC2127,
    _NC2128,
    _NC2129,
    _NC2130,
    _NC2131,
    _NC2132,
    _NC2133,
    _NC2134,
    _NC2135,
    _NC2136,
    _NC2137,
    _NC2138,
    _NC2139,
    _NC2140,
    _NC2141,
    _NC2142,
    _NC2143,
    _NC2144,
    _NC2145,
    _NC2146,
    _NC2147,
    _NC2148,
    _NC2149,
    _NC2150,
    _NC2151,
    _NC2152,
    _NC2153,
    _NC2154,
    _NC2155,
    _NC2156,
    _NC2157,
    _NC2158,
    _NC2159,
    _NC2160,
    _NC2161,
    _NC2162,
    _NC2163,
    _NC2164,
    _NC2165,
    _NC2166}),
    .l15_transducer_data_3({_NC2167,
    _NC2168,
    _NC2169,
    _NC2170,
    _NC2171,
    _NC2172,
    _NC2173,
    _NC2174,
    _NC2175,
    _NC2176,
    _NC2177,
    _NC2178,
    _NC2179,
    _NC2180,
    _NC2181,
    _NC2182,
    _NC2183,
    _NC2184,
    _NC2185,
    _NC2186,
    _NC2187,
    _NC2188,
    _NC2189,
    _NC2190,
    _NC2191,
    _NC2192,
    _NC2193,
    _NC2194,
    _NC2195,
    _NC2196,
    _NC2197,
    _NC2198,
    _NC2199,
    _NC2200,
    _NC2201,
    _NC2202,
    _NC2203,
    _NC2204,
    _NC2205,
    _NC2206,
    _NC2207,
    _NC2208,
    _NC2209,
    _NC2210,
    _NC2211,
    _NC2212,
    _NC2213,
    _NC2214,
    _NC2215,
    _NC2216,
    _NC2217,
    _NC2218,
    _NC2219,
    _NC2220,
    _NC2221,
    _NC2222,
    _NC2223,
    _NC2224,
    _NC2225,
    _NC2226,
    _NC2227,
    _NC2228,
    _NC2229,
    _NC2230}),
    .l15_transducer_error({_NC2231,
    _NC2232}),
    .l15_transducer_inval_address_15_4({_NC2233,
    _NC2234,
    _NC2235,
    _NC2236,
    _NC2237,
    _NC2238,
    _NC2239,
    _NC2240,
    _NC2241,
    _NC2242,
    _NC2243,
    _NC2244}),
    .l15_transducer_inval_way({_NC2245,
    _NC2246}),
    .l15_transducer_returntype({_NC2247,
    _NC2248,
    _NC2249,
    _NC2250}),
    .l2_rtap_data({_NC2251,
    _NC2252,
    _NC2253,
    _NC2254}),
    .noc1_out_data({_NC2255,
    _NC2256,
    _NC2257,
    _NC2258,
    _NC2259,
    _NC2260,
    _NC2261,
    _NC2262,
    _NC2263,
    _NC2264,
    _NC2265,
    _NC2266,
    _NC2267,
    _NC2268,
    _NC2269,
    _NC2270,
    _NC2271,
    _NC2272,
    _NC2273,
    _NC2274,
    _NC2275,
    _NC2276,
    _NC2277,
    _NC2278,
    _NC2279,
    _NC2280,
    _NC2281,
    _NC2282,
    _NC2283,
    _NC2284,
    _NC2285,
    _NC2286,
    _NC2287,
    _NC2288,
    _NC2289,
    _NC2290,
    _NC2291,
    _NC2292,
    _NC2293,
    _NC2294,
    _NC2295,
    _NC2296,
    _NC2297,
    _NC2298,
    _NC2299,
    _NC2300,
    _NC2301,
    _NC2302,
    _NC2303,
    _NC2304,
    _NC2305,
    _NC2306,
    _NC2307,
    _NC2308,
    _NC2309,
    _NC2310,
    _NC2311,
    _NC2312,
    _NC2313,
    _NC2314,
    _NC2315,
    _NC2316,
    _NC2317,
    _NC2318}),
    .noc2_in_data({_NC2319,
    _NC2320,
    _NC2321,
    _NC2322,
    _NC2323,
    _NC2324,
    _NC2325,
    _NC2326,
    _NC2327,
    _NC2328,
    _NC2329,
    _NC2330,
    _NC2331,
    _NC2332,
    _NC2333,
    _NC2334,
    _NC2335,
    _NC2336,
    _NC2337,
    _NC2338,
    _NC2339,
    _NC2340,
    _NC2341,
    _NC2342,
    _NC2343,
    _NC2344,
    _NC2345,
    _NC2346,
    _NC2347,
    _NC2348,
    _NC2349,
    _NC2350,
    _NC2351,
    _NC2352,
    _NC2353,
    _NC2354,
    _NC2355,
    _NC2356,
    _NC2357,
    _NC2358,
    _NC2359,
    _NC2360,
    _NC2361,
    _NC2362,
    _NC2363,
    _NC2364,
    _NC2365,
    _NC2366,
    _NC2367,
    _NC2368,
    _NC2369,
    _NC2370,
    _NC2371,
    _NC2372,
    _NC2373,
    _NC2374,
    _NC2375,
    _NC2376,
    _NC2377,
    _NC2378,
    _NC2379,
    _NC2380,
    _NC2381,
    _NC2382}),
    .noc3_out_data({_NC2383,
    _NC2384,
    _NC2385,
    _NC2386,
    _NC2387,
    _NC2388,
    _NC2389,
    _NC2390,
    _NC2391,
    _NC2392,
    _NC2393,
    _NC2394,
    _NC2395,
    _NC2396,
    _NC2397,
    _NC2398,
    _NC2399,
    _NC2400,
    _NC2401,
    _NC2402,
    _NC2403,
    _NC2404,
    _NC2405,
    _NC2406,
    _NC2407,
    _NC2408,
    _NC2409,
    _NC2410,
    _NC2411,
    _NC2412,
    _NC2413,
    _NC2414,
    _NC2415,
    _NC2416,
    _NC2417,
    _NC2418,
    _NC2419,
    _NC2420,
    _NC2421,
    _NC2422,
    _NC2423,
    _NC2424,
    _NC2425,
    _NC2426,
    _NC2427,
    _NC2428,
    _NC2429,
    _NC2430,
    _NC2431,
    _NC2432,
    _NC2433,
    _NC2434,
    _NC2435,
    _NC2436,
    _NC2437,
    _NC2438,
    _NC2439,
    _NC2440,
    _NC2441,
    _NC2442,
    _NC2443,
    _NC2444,
    _NC2445,
    _NC2446}),
    .processor_router_data_noc2({_NC2447,
    _NC2448,
    _NC2449,
    _NC2450,
    _NC2451,
    _NC2452,
    _NC2453,
    _NC2454,
    _NC2455,
    _NC2456,
    _NC2457,
    _NC2458,
    _NC2459,
    _NC2460,
    _NC2461,
    _NC2462,
    _NC2463,
    _NC2464,
    _NC2465,
    _NC2466,
    _NC2467,
    _NC2468,
    _NC2469,
    _NC2470,
    _NC2471,
    _NC2472,
    _NC2473,
    _NC2474,
    _NC2475,
    _NC2476,
    _NC2477,
    _NC2478,
    _NC2479,
    _NC2480,
    _NC2481,
    _NC2482,
    _NC2483,
    _NC2484,
    _NC2485,
    _NC2486,
    _NC2487,
    _NC2488,
    _NC2489,
    _NC2490,
    _NC2491,
    _NC2492,
    _NC2493,
    _NC2494,
    _NC2495,
    _NC2496,
    _NC2497,
    _NC2498,
    _NC2499,
    _NC2500,
    _NC2501,
    _NC2502,
    _NC2503,
    _NC2504,
    _NC2505,
    _NC2506,
    _NC2507,
    _NC2508,
    _NC2509,
    _NC2510}),
    .rtap_srams_bist_command({_NC2511,
    _NC2512,
    _NC2513,
    _NC2514}),
    .rtap_srams_bist_data({_NC2515,
    _NC2516,
    _NC2517,
    _NC2518}),
    .srams_rtap_data({_NC2519,
    _NC2520,
    _NC2521,
    _NC2522}),
    .tile_jtag_ucb_data({_NC2523,
    _NC2524,
    _NC2525,
    _NC2526}),
    .transducer_l15_address({_NC2527,
    _NC2528,
    _NC2529,
    _NC2530,
    _NC2531,
    _NC2532,
    _NC2533,
    _NC2534,
    _NC2535,
    _NC2536,
    _NC2537,
    _NC2538,
    _NC2539,
    _NC2540,
    _NC2541,
    _NC2542,
    _NC2543,
    _NC2544,
    _NC2545,
    _NC2546,
    _NC2547,
    _NC2548,
    _NC2549,
    _NC2550,
    _NC2551,
    _NC2552,
    _NC2553,
    _NC2554,
    _NC2555,
    _NC2556,
    _NC2557,
    _NC2558,
    _NC2559,
    _NC2560,
    _NC2561,
    _NC2562,
    _NC2563,
    _NC2564,
    _NC2565,
    _NC2566}),
    .transducer_l15_amo_op({_NC2567,
    _NC2568,
    _NC2569,
    _NC2570}),
    .transducer_l15_csm_data({_NC2571,
    _NC2572,
    _NC2573,
    _NC2574,
    _NC2575,
    _NC2576,
    _NC2577,
    _NC2578,
    _NC2579,
    _NC2580,
    _NC2581,
    _NC2582,
    _NC2583,
    _NC2584,
    _NC2585,
    _NC2586,
    _NC2587,
    _NC2588,
    _NC2589,
    _NC2590,
    _NC2591,
    _NC2592,
    _NC2593,
    _NC2594,
    _NC2595,
    _NC2596,
    _NC2597,
    _NC2598,
    _NC2599,
    _NC2600,
    _NC2601,
    _NC2602,
    _NC2603}),
    .transducer_l15_data({_NC2604,
    _NC2605,
    _NC2606,
    _NC2607,
    _NC2608,
    _NC2609,
    _NC2610,
    _NC2611,
    _NC2612,
    _NC2613,
    _NC2614,
    _NC2615,
    _NC2616,
    _NC2617,
    _NC2618,
    _NC2619,
    _NC2620,
    _NC2621,
    _NC2622,
    _NC2623,
    _NC2624,
    _NC2625,
    _NC2626,
    _NC2627,
    _NC2628,
    _NC2629,
    _NC2630,
    _NC2631,
    _NC2632,
    _NC2633,
    _NC2634,
    _NC2635,
    _NC2636,
    _NC2637,
    _NC2638,
    _NC2639,
    _NC2640,
    _NC2641,
    _NC2642,
    _NC2643,
    _NC2644,
    _NC2645,
    _NC2646,
    _NC2647,
    _NC2648,
    _NC2649,
    _NC2650,
    _NC2651,
    _NC2652,
    _NC2653,
    _NC2654,
    _NC2655,
    _NC2656,
    _NC2657,
    _NC2658,
    _NC2659,
    _NC2660,
    _NC2661,
    _NC2662,
    _NC2663,
    _NC2664,
    _NC2665,
    _NC2666,
    _NC2667}),
    .transducer_l15_data_next_entry({_NC2668,
    _NC2669,
    _NC2670,
    _NC2671,
    _NC2672,
    _NC2673,
    _NC2674,
    _NC2675,
    _NC2676,
    _NC2677,
    _NC2678,
    _NC2679,
    _NC2680,
    _NC2681,
    _NC2682,
    _NC2683,
    _NC2684,
    _NC2685,
    _NC2686,
    _NC2687,
    _NC2688,
    _NC2689,
    _NC2690,
    _NC2691,
    _NC2692,
    _NC2693,
    _NC2694,
    _NC2695,
    _NC2696,
    _NC2697,
    _NC2698,
    _NC2699,
    _NC2700,
    _NC2701,
    _NC2702,
    _NC2703,
    _NC2704,
    _NC2705,
    _NC2706,
    _NC2707,
    _NC2708,
    _NC2709,
    _NC2710,
    _NC2711,
    _NC2712,
    _NC2713,
    _NC2714,
    _NC2715,
    _NC2716,
    _NC2717,
    _NC2718,
    _NC2719,
    _NC2720,
    _NC2721,
    _NC2722,
    _NC2723,
    _NC2724,
    _NC2725,
    _NC2726,
    _NC2727,
    _NC2728,
    _NC2729,
    _NC2730,
    _NC2731}),
    .transducer_l15_l1rplway({_NC2732,
    _NC2733}),
    .transducer_l15_rqtype({_NC2734,
    _NC2735,
    _NC2736,
    _NC2737,
    _NC2738}),
    .transducer_l15_size({_NC2739,
    _NC2740,
    _NC2741}));
endmodule

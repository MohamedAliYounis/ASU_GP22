VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tile
  CLASS BLOCK ;
  FOREIGN tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 2500.000 ;
  PIN buffer_processor_data_noc1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 0.000 1919.490 4.000 ;
    END
  END buffer_processor_data_noc1[0]
  PIN buffer_processor_data_noc1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END buffer_processor_data_noc1[10]
  PIN buffer_processor_data_noc1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1009.840 2500.000 1010.440 ;
    END
  END buffer_processor_data_noc1[11]
  PIN buffer_processor_data_noc1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 2496.000 515.570 2500.000 ;
    END
  END buffer_processor_data_noc1[12]
  PIN buffer_processor_data_noc1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1679.640 2500.000 1680.240 ;
    END
  END buffer_processor_data_noc1[13]
  PIN buffer_processor_data_noc1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2352.840 2500.000 2353.440 ;
    END
  END buffer_processor_data_noc1[14]
  PIN buffer_processor_data_noc1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.970 2496.000 1945.250 2500.000 ;
    END
  END buffer_processor_data_noc1[15]
  PIN buffer_processor_data_noc1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 2496.000 837.570 2500.000 ;
    END
  END buffer_processor_data_noc1[16]
  PIN buffer_processor_data_noc1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END buffer_processor_data_noc1[17]
  PIN buffer_processor_data_noc1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 2496.000 1822.890 2500.000 ;
    END
  END buffer_processor_data_noc1[18]
  PIN buffer_processor_data_noc1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.970 2496.000 2428.250 2500.000 ;
    END
  END buffer_processor_data_noc1[19]
  PIN buffer_processor_data_noc1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END buffer_processor_data_noc1[1]
  PIN buffer_processor_data_noc1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END buffer_processor_data_noc1[20]
  PIN buffer_processor_data_noc1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1666.040 2500.000 1666.640 ;
    END
  END buffer_processor_data_noc1[21]
  PIN buffer_processor_data_noc1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2390.240 2500.000 2390.840 ;
    END
  END buffer_processor_data_noc1[22]
  PIN buffer_processor_data_noc1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END buffer_processor_data_noc1[23]
  PIN buffer_processor_data_noc1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2046.840 2500.000 2047.440 ;
    END
  END buffer_processor_data_noc1[24]
  PIN buffer_processor_data_noc1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END buffer_processor_data_noc1[25]
  PIN buffer_processor_data_noc1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 2496.000 225.770 2500.000 ;
    END
  END buffer_processor_data_noc1[26]
  PIN buffer_processor_data_noc1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END buffer_processor_data_noc1[27]
  PIN buffer_processor_data_noc1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END buffer_processor_data_noc1[28]
  PIN buffer_processor_data_noc1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 4.000 ;
    END
  END buffer_processor_data_noc1[29]
  PIN buffer_processor_data_noc1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 0.000 1603.930 4.000 ;
    END
  END buffer_processor_data_noc1[2]
  PIN buffer_processor_data_noc1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1190.040 2500.000 1190.640 ;
    END
  END buffer_processor_data_noc1[30]
  PIN buffer_processor_data_noc1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1540.240 2500.000 1540.840 ;
    END
  END buffer_processor_data_noc1[31]
  PIN buffer_processor_data_noc1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END buffer_processor_data_noc1[32]
  PIN buffer_processor_data_noc1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END buffer_processor_data_noc1[33]
  PIN buffer_processor_data_noc1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 4.000 ;
    END
  END buffer_processor_data_noc1[34]
  PIN buffer_processor_data_noc1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1734.040 4.000 1734.640 ;
    END
  END buffer_processor_data_noc1[35]
  PIN buffer_processor_data_noc1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 2496.000 1053.310 2500.000 ;
    END
  END buffer_processor_data_noc1[36]
  PIN buffer_processor_data_noc1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END buffer_processor_data_noc1[37]
  PIN buffer_processor_data_noc1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END buffer_processor_data_noc1[38]
  PIN buffer_processor_data_noc1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END buffer_processor_data_noc1[39]
  PIN buffer_processor_data_noc1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1584.440 2500.000 1585.040 ;
    END
  END buffer_processor_data_noc1[3]
  PIN buffer_processor_data_noc1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1074.440 2500.000 1075.040 ;
    END
  END buffer_processor_data_noc1[40]
  PIN buffer_processor_data_noc1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 2496.000 161.370 2500.000 ;
    END
  END buffer_processor_data_noc1[41]
  PIN buffer_processor_data_noc1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 0.000 2125.570 4.000 ;
    END
  END buffer_processor_data_noc1[42]
  PIN buffer_processor_data_noc1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1751.040 2500.000 1751.640 ;
    END
  END buffer_processor_data_noc1[43]
  PIN buffer_processor_data_noc1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END buffer_processor_data_noc1[44]
  PIN buffer_processor_data_noc1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END buffer_processor_data_noc1[45]
  PIN buffer_processor_data_noc1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END buffer_processor_data_noc1[46]
  PIN buffer_processor_data_noc1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END buffer_processor_data_noc1[47]
  PIN buffer_processor_data_noc1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 425.040 2500.000 425.640 ;
    END
  END buffer_processor_data_noc1[48]
  PIN buffer_processor_data_noc1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 2496.000 1227.190 2500.000 ;
    END
  END buffer_processor_data_noc1[49]
  PIN buffer_processor_data_noc1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1128.840 2500.000 1129.440 ;
    END
  END buffer_processor_data_noc1[4]
  PIN buffer_processor_data_noc1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2332.440 2500.000 2333.040 ;
    END
  END buffer_processor_data_noc1[50]
  PIN buffer_processor_data_noc1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END buffer_processor_data_noc1[51]
  PIN buffer_processor_data_noc1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 2496.000 2199.630 2500.000 ;
    END
  END buffer_processor_data_noc1[52]
  PIN buffer_processor_data_noc1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END buffer_processor_data_noc1[53]
  PIN buffer_processor_data_noc1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END buffer_processor_data_noc1[54]
  PIN buffer_processor_data_noc1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 2496.000 280.510 2500.000 ;
    END
  END buffer_processor_data_noc1[55]
  PIN buffer_processor_data_noc1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1870.040 2500.000 1870.640 ;
    END
  END buffer_processor_data_noc1[56]
  PIN buffer_processor_data_noc1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END buffer_processor_data_noc1[57]
  PIN buffer_processor_data_noc1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END buffer_processor_data_noc1[58]
  PIN buffer_processor_data_noc1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 2496.000 1742.390 2500.000 ;
    END
  END buffer_processor_data_noc1[59]
  PIN buffer_processor_data_noc1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.330 0.000 2067.610 4.000 ;
    END
  END buffer_processor_data_noc1[5]
  PIN buffer_processor_data_noc1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END buffer_processor_data_noc1[60]
  PIN buffer_processor_data_noc1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 0.000 1259.390 4.000 ;
    END
  END buffer_processor_data_noc1[61]
  PIN buffer_processor_data_noc1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.710 2496.000 1838.990 2500.000 ;
    END
  END buffer_processor_data_noc1[62]
  PIN buffer_processor_data_noc1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END buffer_processor_data_noc1[63]
  PIN buffer_processor_data_noc1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.990 0.000 2399.270 4.000 ;
    END
  END buffer_processor_data_noc1[6]
  PIN buffer_processor_data_noc1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END buffer_processor_data_noc1[7]
  PIN buffer_processor_data_noc1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 2496.000 979.250 2500.000 ;
    END
  END buffer_processor_data_noc1[8]
  PIN buffer_processor_data_noc1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 2496.000 1143.470 2500.000 ;
    END
  END buffer_processor_data_noc1[9]
  PIN buffer_processor_data_noc3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END buffer_processor_data_noc3[0]
  PIN buffer_processor_data_noc3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2254.240 2500.000 2254.840 ;
    END
  END buffer_processor_data_noc3[10]
  PIN buffer_processor_data_noc3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 799.040 2500.000 799.640 ;
    END
  END buffer_processor_data_noc3[11]
  PIN buffer_processor_data_noc3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 2496.000 1694.090 2500.000 ;
    END
  END buffer_processor_data_noc3[12]
  PIN buffer_processor_data_noc3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 2496.000 67.990 2500.000 ;
    END
  END buffer_processor_data_noc3[13]
  PIN buffer_processor_data_noc3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 44.240 2500.000 44.840 ;
    END
  END buffer_processor_data_noc3[14]
  PIN buffer_processor_data_noc3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 2496.000 1291.590 2500.000 ;
    END
  END buffer_processor_data_noc3[15]
  PIN buffer_processor_data_noc3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.590 2496.000 2173.870 2500.000 ;
    END
  END buffer_processor_data_noc3[16]
  PIN buffer_processor_data_noc3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END buffer_processor_data_noc3[17]
  PIN buffer_processor_data_noc3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1604.840 2500.000 1605.440 ;
    END
  END buffer_processor_data_noc3[18]
  PIN buffer_processor_data_noc3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.770 0.000 2074.050 4.000 ;
    END
  END buffer_processor_data_noc3[19]
  PIN buffer_processor_data_noc3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 445.440 2500.000 446.040 ;
    END
  END buffer_processor_data_noc3[1]
  PIN buffer_processor_data_noc3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END buffer_processor_data_noc3[20]
  PIN buffer_processor_data_noc3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2186.240 4.000 2186.840 ;
    END
  END buffer_processor_data_noc3[21]
  PIN buffer_processor_data_noc3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1951.640 2500.000 1952.240 ;
    END
  END buffer_processor_data_noc3[22]
  PIN buffer_processor_data_noc3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1812.240 4.000 1812.840 ;
    END
  END buffer_processor_data_noc3[23]
  PIN buffer_processor_data_noc3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2203.240 4.000 2203.840 ;
    END
  END buffer_processor_data_noc3[24]
  PIN buffer_processor_data_noc3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 867.040 2500.000 867.640 ;
    END
  END buffer_processor_data_noc3[25]
  PIN buffer_processor_data_noc3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 0.000 1568.510 4.000 ;
    END
  END buffer_processor_data_noc3[26]
  PIN buffer_processor_data_noc3[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END buffer_processor_data_noc3[27]
  PIN buffer_processor_data_noc3[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 748.040 2500.000 748.640 ;
    END
  END buffer_processor_data_noc3[28]
  PIN buffer_processor_data_noc3[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END buffer_processor_data_noc3[29]
  PIN buffer_processor_data_noc3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1662.640 4.000 1663.240 ;
    END
  END buffer_processor_data_noc3[2]
  PIN buffer_processor_data_noc3[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END buffer_processor_data_noc3[30]
  PIN buffer_processor_data_noc3[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END buffer_processor_data_noc3[31]
  PIN buffer_processor_data_noc3[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END buffer_processor_data_noc3[32]
  PIN buffer_processor_data_noc3[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 0.000 1188.550 4.000 ;
    END
  END buffer_processor_data_noc3[33]
  PIN buffer_processor_data_noc3[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END buffer_processor_data_noc3[34]
  PIN buffer_processor_data_noc3[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 809.240 2500.000 809.840 ;
    END
  END buffer_processor_data_noc3[35]
  PIN buffer_processor_data_noc3[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 880.640 2500.000 881.240 ;
    END
  END buffer_processor_data_noc3[36]
  PIN buffer_processor_data_noc3[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1822.440 2500.000 1823.040 ;
    END
  END buffer_processor_data_noc3[37]
  PIN buffer_processor_data_noc3[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END buffer_processor_data_noc3[38]
  PIN buffer_processor_data_noc3[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.030 0.000 2180.310 4.000 ;
    END
  END buffer_processor_data_noc3[39]
  PIN buffer_processor_data_noc3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.870 0.000 2251.150 4.000 ;
    END
  END buffer_processor_data_noc3[3]
  PIN buffer_processor_data_noc3[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 2496.000 1407.510 2500.000 ;
    END
  END buffer_processor_data_noc3[40]
  PIN buffer_processor_data_noc3[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END buffer_processor_data_noc3[41]
  PIN buffer_processor_data_noc3[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 2496.000 1568.510 2500.000 ;
    END
  END buffer_processor_data_noc3[42]
  PIN buffer_processor_data_noc3[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 0.000 2012.870 4.000 ;
    END
  END buffer_processor_data_noc3[43]
  PIN buffer_processor_data_noc3[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 414.840 2500.000 415.440 ;
    END
  END buffer_processor_data_noc3[44]
  PIN buffer_processor_data_noc3[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1720.440 2500.000 1721.040 ;
    END
  END buffer_processor_data_noc3[45]
  PIN buffer_processor_data_noc3[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 0.000 1942.030 4.000 ;
    END
  END buffer_processor_data_noc3[46]
  PIN buffer_processor_data_noc3[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END buffer_processor_data_noc3[47]
  PIN buffer_processor_data_noc3[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END buffer_processor_data_noc3[48]
  PIN buffer_processor_data_noc3[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.290 0.000 1803.570 4.000 ;
    END
  END buffer_processor_data_noc3[49]
  PIN buffer_processor_data_noc3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 2496.000 596.070 2500.000 ;
    END
  END buffer_processor_data_noc3[4]
  PIN buffer_processor_data_noc3[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END buffer_processor_data_noc3[50]
  PIN buffer_processor_data_noc3[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2148.840 4.000 2149.440 ;
    END
  END buffer_processor_data_noc3[51]
  PIN buffer_processor_data_noc3[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END buffer_processor_data_noc3[52]
  PIN buffer_processor_data_noc3[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 4.000 ;
    END
  END buffer_processor_data_noc3[53]
  PIN buffer_processor_data_noc3[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1706.840 4.000 1707.440 ;
    END
  END buffer_processor_data_noc3[54]
  PIN buffer_processor_data_noc3[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END buffer_processor_data_noc3[55]
  PIN buffer_processor_data_noc3[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END buffer_processor_data_noc3[56]
  PIN buffer_processor_data_noc3[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 0.000 1037.210 4.000 ;
    END
  END buffer_processor_data_noc3[57]
  PIN buffer_processor_data_noc3[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END buffer_processor_data_noc3[58]
  PIN buffer_processor_data_noc3[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END buffer_processor_data_noc3[59]
  PIN buffer_processor_data_noc3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1098.240 2500.000 1098.840 ;
    END
  END buffer_processor_data_noc3[5]
  PIN buffer_processor_data_noc3[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END buffer_processor_data_noc3[60]
  PIN buffer_processor_data_noc3[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.270 2496.000 1993.550 2500.000 ;
    END
  END buffer_processor_data_noc3[61]
  PIN buffer_processor_data_noc3[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END buffer_processor_data_noc3[62]
  PIN buffer_processor_data_noc3[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 2496.000 42.230 2500.000 ;
    END
  END buffer_processor_data_noc3[63]
  PIN buffer_processor_data_noc3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END buffer_processor_data_noc3[6]
  PIN buffer_processor_data_noc3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END buffer_processor_data_noc3[7]
  PIN buffer_processor_data_noc3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END buffer_processor_data_noc3[8]
  PIN buffer_processor_data_noc3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 2496.000 2135.230 2500.000 ;
    END
  END buffer_processor_data_noc3[9]
  PIN buffer_processor_valid_noc1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 71.440 2500.000 72.040 ;
    END
  END buffer_processor_valid_noc1
  PIN buffer_processor_valid_noc3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END buffer_processor_valid_noc3
  PIN chipid[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.240 4.000 1438.840 ;
    END
  END chipid[0]
  PIN chipid[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END chipid[10]
  PIN chipid[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 0.000 1516.990 4.000 ;
    END
  END chipid[11]
  PIN chipid[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END chipid[12]
  PIN chipid[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END chipid[13]
  PIN chipid[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END chipid[1]
  PIN chipid[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.410 2496.000 1951.690 2500.000 ;
    END
  END chipid[2]
  PIN chipid[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2050.240 4.000 2050.840 ;
    END
  END chipid[3]
  PIN chipid[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END chipid[4]
  PIN chipid[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END chipid[5]
  PIN chipid[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.390 0.000 1819.670 4.000 ;
    END
  END chipid[6]
  PIN chipid[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 2496.000 1954.910 2500.000 ;
    END
  END chipid[7]
  PIN chipid[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2469.830 0.000 2470.110 4.000 ;
    END
  END chipid[8]
  PIN chipid[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 2496.000 992.130 2500.000 ;
    END
  END chipid[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 238.040 2500.000 238.640 ;
    END
  END clk
  PIN clk_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 2496.000 1352.770 2500.000 ;
    END
  END clk_en
  PIN config_chipid[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END config_chipid[0]
  PIN config_chipid[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 2496.000 1584.610 2500.000 ;
    END
  END config_chipid[10]
  PIN config_chipid[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END config_chipid[11]
  PIN config_chipid[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END config_chipid[12]
  PIN config_chipid[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 887.440 2500.000 888.040 ;
    END
  END config_chipid[13]
  PIN config_chipid[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 2496.000 1314.130 2500.000 ;
    END
  END config_chipid[1]
  PIN config_chipid[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 2496.000 1030.770 2500.000 ;
    END
  END config_chipid[2]
  PIN config_chipid[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END config_chipid[3]
  PIN config_chipid[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END config_chipid[4]
  PIN config_chipid[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 2496.000 1104.830 2500.000 ;
    END
  END config_chipid[5]
  PIN config_chipid[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 0.000 1790.690 4.000 ;
    END
  END config_chipid[6]
  PIN config_chipid[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 4.000 ;
    END
  END config_chipid[7]
  PIN config_chipid[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 2496.000 2160.990 2500.000 ;
    END
  END config_chipid[8]
  PIN config_chipid[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1982.240 4.000 1982.840 ;
    END
  END config_chipid[9]
  PIN config_coreid_x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 289.040 2500.000 289.640 ;
    END
  END config_coreid_x[0]
  PIN config_coreid_x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1084.640 2500.000 1085.240 ;
    END
  END config_coreid_x[1]
  PIN config_coreid_x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.630 0.000 2437.910 4.000 ;
    END
  END config_coreid_x[2]
  PIN config_coreid_x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 0.000 2160.990 4.000 ;
    END
  END config_coreid_x[3]
  PIN config_coreid_x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2135.240 2500.000 2135.840 ;
    END
  END config_coreid_x[4]
  PIN config_coreid_x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END config_coreid_x[5]
  PIN config_coreid_x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1526.640 4.000 1527.240 ;
    END
  END config_coreid_x[6]
  PIN config_coreid_x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END config_coreid_x[7]
  PIN config_coreid_y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 2496.000 969.590 2500.000 ;
    END
  END config_coreid_y[0]
  PIN config_coreid_y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END config_coreid_y[1]
  PIN config_coreid_y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 2496.000 625.050 2500.000 ;
    END
  END config_coreid_y[2]
  PIN config_coreid_y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END config_coreid_y[3]
  PIN config_coreid_y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END config_coreid_y[4]
  PIN config_coreid_y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END config_coreid_y[5]
  PIN config_coreid_y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 649.440 2500.000 650.040 ;
    END
  END config_coreid_y[6]
  PIN config_coreid_y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1791.840 2500.000 1792.440 ;
    END
  END config_coreid_y[7]
  PIN config_csm_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2189.640 2500.000 2190.240 ;
    END
  END config_csm_en
  PIN config_hmt_base[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690 2496.000 2350.970 2500.000 ;
    END
  END config_hmt_base[0]
  PIN config_hmt_base[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END config_hmt_base[10]
  PIN config_hmt_base[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.370 2496.000 2009.650 2500.000 ;
    END
  END config_hmt_base[11]
  PIN config_hmt_base[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 0.000 2225.390 4.000 ;
    END
  END config_hmt_base[12]
  PIN config_hmt_base[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1951.640 4.000 1952.240 ;
    END
  END config_hmt_base[13]
  PIN config_hmt_base[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 2496.000 1288.370 2500.000 ;
    END
  END config_hmt_base[14]
  PIN config_hmt_base[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 2496.000 10.030 2500.000 ;
    END
  END config_hmt_base[15]
  PIN config_hmt_base[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END config_hmt_base[16]
  PIN config_hmt_base[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1567.440 2500.000 1568.040 ;
    END
  END config_hmt_base[17]
  PIN config_hmt_base[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 2496.000 1797.130 2500.000 ;
    END
  END config_hmt_base[18]
  PIN config_hmt_base[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 2496.000 486.590 2500.000 ;
    END
  END config_hmt_base[19]
  PIN config_hmt_base[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2162.440 4.000 2163.040 ;
    END
  END config_hmt_base[1]
  PIN config_hmt_base[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END config_hmt_base[20]
  PIN config_hmt_base[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 2496.000 109.850 2500.000 ;
    END
  END config_hmt_base[21]
  PIN config_hmt_base[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 2496.000 74.430 2500.000 ;
    END
  END config_hmt_base[2]
  PIN config_hmt_base[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 2496.000 1317.350 2500.000 ;
    END
  END config_hmt_base[3]
  PIN config_hmt_base[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 0.000 1339.890 4.000 ;
    END
  END config_hmt_base[4]
  PIN config_hmt_base[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 2496.000 1198.210 2500.000 ;
    END
  END config_hmt_base[5]
  PIN config_hmt_base[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END config_hmt_base[6]
  PIN config_hmt_base[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 472.640 2500.000 473.240 ;
    END
  END config_hmt_base[7]
  PIN config_hmt_base[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 2496.000 1037.210 2500.000 ;
    END
  END config_hmt_base[8]
  PIN config_hmt_base[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END config_hmt_base[9]
  PIN config_home_alloc_method[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END config_home_alloc_method[0]
  PIN config_home_alloc_method[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1118.640 2500.000 1119.240 ;
    END
  END config_home_alloc_method[1]
  PIN config_l15_read_res_data_s3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 2496.000 1182.110 2500.000 ;
    END
  END config_l15_read_res_data_s3[0]
  PIN config_l15_read_res_data_s3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.590 2496.000 2334.870 2500.000 ;
    END
  END config_l15_read_res_data_s3[10]
  PIN config_l15_read_res_data_s3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 2496.000 422.190 2500.000 ;
    END
  END config_l15_read_res_data_s3[11]
  PIN config_l15_read_res_data_s3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1819.040 2500.000 1819.640 ;
    END
  END config_l15_read_res_data_s3[12]
  PIN config_l15_read_res_data_s3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2397.040 2500.000 2397.640 ;
    END
  END config_l15_read_res_data_s3[13]
  PIN config_l15_read_res_data_s3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 340.040 2500.000 340.640 ;
    END
  END config_l15_read_res_data_s3[14]
  PIN config_l15_read_res_data_s3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 2496.000 55.110 2500.000 ;
    END
  END config_l15_read_res_data_s3[15]
  PIN config_l15_read_res_data_s3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 2496.000 1507.330 2500.000 ;
    END
  END config_l15_read_res_data_s3[16]
  PIN config_l15_read_res_data_s3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 2496.000 219.330 2500.000 ;
    END
  END config_l15_read_res_data_s3[17]
  PIN config_l15_read_res_data_s3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END config_l15_read_res_data_s3[18]
  PIN config_l15_read_res_data_s3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END config_l15_read_res_data_s3[19]
  PIN config_l15_read_res_data_s3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END config_l15_read_res_data_s3[1]
  PIN config_l15_read_res_data_s3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END config_l15_read_res_data_s3[20]
  PIN config_l15_read_res_data_s3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END config_l15_read_res_data_s3[21]
  PIN config_l15_read_res_data_s3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END config_l15_read_res_data_s3[22]
  PIN config_l15_read_res_data_s3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1659.240 4.000 1659.840 ;
    END
  END config_l15_read_res_data_s3[23]
  PIN config_l15_read_res_data_s3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2165.840 2500.000 2166.440 ;
    END
  END config_l15_read_res_data_s3[24]
  PIN config_l15_read_res_data_s3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1836.040 2500.000 1836.640 ;
    END
  END config_l15_read_res_data_s3[25]
  PIN config_l15_read_res_data_s3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.930 2496.000 2164.210 2500.000 ;
    END
  END config_l15_read_res_data_s3[26]
  PIN config_l15_read_res_data_s3[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END config_l15_read_res_data_s3[27]
  PIN config_l15_read_res_data_s3[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 0.000 1423.610 4.000 ;
    END
  END config_l15_read_res_data_s3[28]
  PIN config_l15_read_res_data_s3[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.040 4.000 1649.640 ;
    END
  END config_l15_read_res_data_s3[29]
  PIN config_l15_read_res_data_s3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2080.840 4.000 2081.440 ;
    END
  END config_l15_read_res_data_s3[2]
  PIN config_l15_read_res_data_s3[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.950 0.000 2296.230 4.000 ;
    END
  END config_l15_read_res_data_s3[30]
  PIN config_l15_read_res_data_s3[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1268.240 2500.000 1268.840 ;
    END
  END config_l15_read_res_data_s3[31]
  PIN config_l15_read_res_data_s3[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 234.640 2500.000 235.240 ;
    END
  END config_l15_read_res_data_s3[32]
  PIN config_l15_read_res_data_s3[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 0.000 1697.310 4.000 ;
    END
  END config_l15_read_res_data_s3[33]
  PIN config_l15_read_res_data_s3[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 2496.000 1684.430 2500.000 ;
    END
  END config_l15_read_res_data_s3[34]
  PIN config_l15_read_res_data_s3[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.370 2496.000 2492.650 2500.000 ;
    END
  END config_l15_read_res_data_s3[35]
  PIN config_l15_read_res_data_s3[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1247.840 2500.000 1248.440 ;
    END
  END config_l15_read_res_data_s3[36]
  PIN config_l15_read_res_data_s3[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END config_l15_read_res_data_s3[37]
  PIN config_l15_read_res_data_s3[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.490 2496.000 2318.770 2500.000 ;
    END
  END config_l15_read_res_data_s3[38]
  PIN config_l15_read_res_data_s3[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END config_l15_read_res_data_s3[39]
  PIN config_l15_read_res_data_s3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 2496.000 13.250 2500.000 ;
    END
  END config_l15_read_res_data_s3[3]
  PIN config_l15_read_res_data_s3[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END config_l15_read_res_data_s3[40]
  PIN config_l15_read_res_data_s3[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 2496.000 277.290 2500.000 ;
    END
  END config_l15_read_res_data_s3[41]
  PIN config_l15_read_res_data_s3[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 955.440 2500.000 956.040 ;
    END
  END config_l15_read_res_data_s3[42]
  PIN config_l15_read_res_data_s3[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 2496.000 1735.950 2500.000 ;
    END
  END config_l15_read_res_data_s3[43]
  PIN config_l15_read_res_data_s3[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 2496.000 1861.530 2500.000 ;
    END
  END config_l15_read_res_data_s3[44]
  PIN config_l15_read_res_data_s3[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 2496.000 1687.650 2500.000 ;
    END
  END config_l15_read_res_data_s3[45]
  PIN config_l15_read_res_data_s3[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END config_l15_read_res_data_s3[46]
  PIN config_l15_read_res_data_s3[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END config_l15_read_res_data_s3[47]
  PIN config_l15_read_res_data_s3[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END config_l15_read_res_data_s3[48]
  PIN config_l15_read_res_data_s3[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 0.000 2080.490 4.000 ;
    END
  END config_l15_read_res_data_s3[49]
  PIN config_l15_read_res_data_s3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 108.840 2500.000 109.440 ;
    END
  END config_l15_read_res_data_s3[4]
  PIN config_l15_read_res_data_s3[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1917.640 4.000 1918.240 ;
    END
  END config_l15_read_res_data_s3[50]
  PIN config_l15_read_res_data_s3[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 2496.000 1323.790 2500.000 ;
    END
  END config_l15_read_res_data_s3[51]
  PIN config_l15_read_res_data_s3[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 2496.000 869.770 2500.000 ;
    END
  END config_l15_read_res_data_s3[52]
  PIN config_l15_read_res_data_s3[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END config_l15_read_res_data_s3[53]
  PIN config_l15_read_res_data_s3[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.930 2496.000 2325.210 2500.000 ;
    END
  END config_l15_read_res_data_s3[54]
  PIN config_l15_read_res_data_s3[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END config_l15_read_res_data_s3[55]
  PIN config_l15_read_res_data_s3[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 0.000 2138.450 4.000 ;
    END
  END config_l15_read_res_data_s3[56]
  PIN config_l15_read_res_data_s3[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END config_l15_read_res_data_s3[57]
  PIN config_l15_read_res_data_s3[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2383.440 4.000 2384.040 ;
    END
  END config_l15_read_res_data_s3[58]
  PIN config_l15_read_res_data_s3[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END config_l15_read_res_data_s3[59]
  PIN config_l15_read_res_data_s3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END config_l15_read_res_data_s3[5]
  PIN config_l15_read_res_data_s3[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END config_l15_read_res_data_s3[60]
  PIN config_l15_read_res_data_s3[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 897.640 2500.000 898.240 ;
    END
  END config_l15_read_res_data_s3[61]
  PIN config_l15_read_res_data_s3[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 571.240 2500.000 571.840 ;
    END
  END config_l15_read_res_data_s3[62]
  PIN config_l15_read_res_data_s3[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 98.640 2500.000 99.240 ;
    END
  END config_l15_read_res_data_s3[63]
  PIN config_l15_read_res_data_s3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END config_l15_read_res_data_s3[6]
  PIN config_l15_read_res_data_s3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1982.240 2500.000 1982.840 ;
    END
  END config_l15_read_res_data_s3[7]
  PIN config_l15_read_res_data_s3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.790 0.000 2206.070 4.000 ;
    END
  END config_l15_read_res_data_s3[8]
  PIN config_l15_read_res_data_s3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END config_l15_read_res_data_s3[9]
  PIN config_system_tile_count_5_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.130 0.000 2196.410 4.000 ;
    END
  END config_system_tile_count_5_0[0]
  PIN config_system_tile_count_5_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END config_system_tile_count_5_0[1]
  PIN config_system_tile_count_5_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 431.840 2500.000 432.440 ;
    END
  END config_system_tile_count_5_0[2]
  PIN config_system_tile_count_5_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END config_system_tile_count_5_0[3]
  PIN config_system_tile_count_5_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END config_system_tile_count_5_0[4]
  PIN config_system_tile_count_5_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 2496.000 35.790 2500.000 ;
    END
  END config_system_tile_count_5_0[5]
  PIN coreid_x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 0.000 1314.130 4.000 ;
    END
  END coreid_x[0]
  PIN coreid_x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1805.440 2500.000 1806.040 ;
    END
  END coreid_x[1]
  PIN coreid_x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 68.040 2500.000 68.640 ;
    END
  END coreid_x[2]
  PIN coreid_x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 2496.000 2186.750 2500.000 ;
    END
  END coreid_x[3]
  PIN coreid_x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1516.440 2500.000 1517.040 ;
    END
  END coreid_x[4]
  PIN coreid_x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 2496.000 1465.470 2500.000 ;
    END
  END coreid_x[5]
  PIN coreid_x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1615.040 4.000 1615.640 ;
    END
  END coreid_x[6]
  PIN coreid_x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1679.640 4.000 1680.240 ;
    END
  END coreid_x[7]
  PIN coreid_y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2159.040 2500.000 2159.640 ;
    END
  END coreid_y[0]
  PIN coreid_y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2482.040 2500.000 2482.640 ;
    END
  END coreid_y[1]
  PIN coreid_y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 204.040 2500.000 204.640 ;
    END
  END coreid_y[2]
  PIN coreid_y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1975.440 2500.000 1976.040 ;
    END
  END coreid_y[3]
  PIN coreid_y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2104.640 4.000 2105.240 ;
    END
  END coreid_y[4]
  PIN coreid_y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1961.840 2500.000 1962.440 ;
    END
  END coreid_y[5]
  PIN coreid_y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 2496.000 22.910 2500.000 ;
    END
  END coreid_y[6]
  PIN coreid_y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1244.440 2500.000 1245.040 ;
    END
  END coreid_y[7]
  PIN default_chipid[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END default_chipid[0]
  PIN default_chipid[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 612.040 2500.000 612.640 ;
    END
  END default_chipid[10]
  PIN default_chipid[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 2496.000 811.810 2500.000 ;
    END
  END default_chipid[11]
  PIN default_chipid[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 2496.000 58.330 2500.000 ;
    END
  END default_chipid[12]
  PIN default_chipid[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 2496.000 1336.670 2500.000 ;
    END
  END default_chipid[13]
  PIN default_chipid[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END default_chipid[1]
  PIN default_chipid[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 901.040 2500.000 901.640 ;
    END
  END default_chipid[2]
  PIN default_chipid[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.040 4.000 1751.640 ;
    END
  END default_chipid[3]
  PIN default_chipid[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END default_chipid[4]
  PIN default_chipid[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2366.440 2500.000 2367.040 ;
    END
  END default_chipid[5]
  PIN default_chipid[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 2496.000 367.450 2500.000 ;
    END
  END default_chipid[6]
  PIN default_chipid[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 2496.000 1298.030 2500.000 ;
    END
  END default_chipid[7]
  PIN default_chipid[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 2496.000 1810.010 2500.000 ;
    END
  END default_chipid[8]
  PIN default_chipid[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1319.240 2500.000 1319.840 ;
    END
  END default_chipid[9]
  PIN default_coreid_x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.310 2496.000 1774.590 2500.000 ;
    END
  END default_coreid_x[0]
  PIN default_coreid_x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END default_coreid_x[1]
  PIN default_coreid_x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END default_coreid_x[2]
  PIN default_coreid_x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 2496.000 1272.270 2500.000 ;
    END
  END default_coreid_x[3]
  PIN default_coreid_x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1907.440 2500.000 1908.040 ;
    END
  END default_coreid_x[4]
  PIN default_coreid_x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END default_coreid_x[5]
  PIN default_coreid_x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 2496.000 2177.090 2500.000 ;
    END
  END default_coreid_x[6]
  PIN default_coreid_x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END default_coreid_x[7]
  PIN default_coreid_y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2193.040 2500.000 2193.640 ;
    END
  END default_coreid_y[0]
  PIN default_coreid_y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1686.440 2500.000 1687.040 ;
    END
  END default_coreid_y[1]
  PIN default_coreid_y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END default_coreid_y[2]
  PIN default_coreid_y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END default_coreid_y[3]
  PIN default_coreid_y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 765.040 2500.000 765.640 ;
    END
  END default_coreid_y[4]
  PIN default_coreid_y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 78.240 2500.000 78.840 ;
    END
  END default_coreid_y[5]
  PIN default_coreid_y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END default_coreid_y[6]
  PIN default_coreid_y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 2496.000 0.370 2500.000 ;
    END
  END default_coreid_y[7]
  PIN dmbr_l15_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 4.000 ;
    END
  END dmbr_l15_stall
  PIN dummy_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 761.640 2500.000 762.240 ;
    END
  END dummy_core[0]
  PIN dummy_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 0.000 1533.090 4.000 ;
    END
  END dummy_core[10]
  PIN dummy_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 0.000 1652.230 4.000 ;
    END
  END dummy_core[11]
  PIN dummy_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END dummy_core[12]
  PIN dummy_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 0.000 1745.610 4.000 ;
    END
  END dummy_core[13]
  PIN dummy_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2026.440 2500.000 2027.040 ;
    END
  END dummy_core[14]
  PIN dummy_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 2496.000 531.670 2500.000 ;
    END
  END dummy_core[15]
  PIN dummy_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END dummy_core[16]
  PIN dummy_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 0.000 1594.270 4.000 ;
    END
  END dummy_core[17]
  PIN dummy_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1611.640 4.000 1612.240 ;
    END
  END dummy_core[18]
  PIN dummy_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2128.440 2500.000 2129.040 ;
    END
  END dummy_core[19]
  PIN dummy_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END dummy_core[1]
  PIN dummy_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.690 2496.000 1384.970 2500.000 ;
    END
  END dummy_core[20]
  PIN dummy_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.930 0.000 2486.210 4.000 ;
    END
  END dummy_core[21]
  PIN dummy_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END dummy_core[22]
  PIN dummy_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END dummy_core[23]
  PIN dummy_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END dummy_core[24]
  PIN dummy_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END dummy_core[25]
  PIN dummy_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.950 2496.000 2457.230 2500.000 ;
    END
  END dummy_core[26]
  PIN dummy_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 2496.000 1806.790 2500.000 ;
    END
  END dummy_core[27]
  PIN dummy_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 965.640 2500.000 966.240 ;
    END
  END dummy_core[28]
  PIN dummy_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2244.040 2500.000 2244.640 ;
    END
  END dummy_core[29]
  PIN dummy_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 833.040 2500.000 833.640 ;
    END
  END dummy_core[2]
  PIN dummy_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.750 0.000 2425.030 4.000 ;
    END
  END dummy_core[30]
  PIN dummy_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 788.840 2500.000 789.440 ;
    END
  END dummy_core[31]
  PIN dummy_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 554.240 2500.000 554.840 ;
    END
  END dummy_core[3]
  PIN dummy_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1305.640 2500.000 1306.240 ;
    END
  END dummy_core[4]
  PIN dummy_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 989.440 4.000 990.040 ;
    END
  END dummy_core[5]
  PIN dummy_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2495.590 0.000 2495.870 4.000 ;
    END
  END dummy_core[6]
  PIN dummy_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1866.640 4.000 1867.240 ;
    END
  END dummy_core[7]
  PIN dummy_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 4.000 ;
    END
  END dummy_core[8]
  PIN dummy_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END dummy_core[9]
  PIN dyn0_dEo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 2496.000 1368.870 2500.000 ;
    END
  END dyn0_dEo[0]
  PIN dyn0_dEo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 669.840 2500.000 670.440 ;
    END
  END dyn0_dEo[10]
  PIN dyn0_dEo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END dyn0_dEo[11]
  PIN dyn0_dEo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1723.840 2500.000 1724.440 ;
    END
  END dyn0_dEo[12]
  PIN dyn0_dEo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 2496.000 26.130 2500.000 ;
    END
  END dyn0_dEo[13]
  PIN dyn0_dEo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END dyn0_dEo[14]
  PIN dyn0_dEo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 380.840 2500.000 381.440 ;
    END
  END dyn0_dEo[15]
  PIN dyn0_dEo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.350 2496.000 1877.630 2500.000 ;
    END
  END dyn0_dEo[16]
  PIN dyn0_dEo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END dyn0_dEo[17]
  PIN dyn0_dEo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1717.040 4.000 1717.640 ;
    END
  END dyn0_dEo[18]
  PIN dyn0_dEo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 0.000 1436.490 4.000 ;
    END
  END dyn0_dEo[19]
  PIN dyn0_dEo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.330 2496.000 2389.610 2500.000 ;
    END
  END dyn0_dEo[1]
  PIN dyn0_dEo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2278.040 2500.000 2278.640 ;
    END
  END dyn0_dEo[20]
  PIN dyn0_dEo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 2496.000 1017.890 2500.000 ;
    END
  END dyn0_dEo[21]
  PIN dyn0_dEo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 2496.000 782.830 2500.000 ;
    END
  END dyn0_dEo[22]
  PIN dyn0_dEo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 2496.000 1262.610 2500.000 ;
    END
  END dyn0_dEo[23]
  PIN dyn0_dEo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 2496.000 312.710 2500.000 ;
    END
  END dyn0_dEo[24]
  PIN dyn0_dEo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 81.640 2500.000 82.240 ;
    END
  END dyn0_dEo[25]
  PIN dyn0_dEo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 0.000 2135.230 4.000 ;
    END
  END dyn0_dEo[26]
  PIN dyn0_dEo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 2496.000 370.670 2500.000 ;
    END
  END dyn0_dEo[27]
  PIN dyn0_dEo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.010 2496.000 2370.290 2500.000 ;
    END
  END dyn0_dEo[28]
  PIN dyn0_dEo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END dyn0_dEo[29]
  PIN dyn0_dEo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END dyn0_dEo[2]
  PIN dyn0_dEo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.710 0.000 1838.990 4.000 ;
    END
  END dyn0_dEo[30]
  PIN dyn0_dEo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1030.240 2500.000 1030.840 ;
    END
  END dyn0_dEo[31]
  PIN dyn0_dEo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 2496.000 264.410 2500.000 ;
    END
  END dyn0_dEo[32]
  PIN dyn0_dEo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 2496.000 71.210 2500.000 ;
    END
  END dyn0_dEo[33]
  PIN dyn0_dEo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END dyn0_dEo[34]
  PIN dyn0_dEo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END dyn0_dEo[35]
  PIN dyn0_dEo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 2496.000 1777.810 2500.000 ;
    END
  END dyn0_dEo[36]
  PIN dyn0_dEo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2329.040 2500.000 2329.640 ;
    END
  END dyn0_dEo[37]
  PIN dyn0_dEo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END dyn0_dEo[38]
  PIN dyn0_dEo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END dyn0_dEo[39]
  PIN dyn0_dEo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END dyn0_dEo[3]
  PIN dyn0_dEo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END dyn0_dEo[40]
  PIN dyn0_dEo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 2496.000 1024.330 2500.000 ;
    END
  END dyn0_dEo[41]
  PIN dyn0_dEo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END dyn0_dEo[42]
  PIN dyn0_dEo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END dyn0_dEo[43]
  PIN dyn0_dEo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 2496.000 892.310 2500.000 ;
    END
  END dyn0_dEo[44]
  PIN dyn0_dEo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 0.000 1842.210 4.000 ;
    END
  END dyn0_dEo[45]
  PIN dyn0_dEo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2414.040 2500.000 2414.640 ;
    END
  END dyn0_dEo[46]
  PIN dyn0_dEo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 2496.000 2070.830 2500.000 ;
    END
  END dyn0_dEo[47]
  PIN dyn0_dEo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2366.790 0.000 2367.070 4.000 ;
    END
  END dyn0_dEo[48]
  PIN dyn0_dEo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 217.640 2500.000 218.240 ;
    END
  END dyn0_dEo[49]
  PIN dyn0_dEo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1604.840 4.000 1605.440 ;
    END
  END dyn0_dEo[4]
  PIN dyn0_dEo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END dyn0_dEo[50]
  PIN dyn0_dEo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.610 0.000 2466.890 4.000 ;
    END
  END dyn0_dEo[51]
  PIN dyn0_dEo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END dyn0_dEo[52]
  PIN dyn0_dEo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END dyn0_dEo[53]
  PIN dyn0_dEo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 2496.000 1426.830 2500.000 ;
    END
  END dyn0_dEo[54]
  PIN dyn0_dEo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 2496.000 605.730 2500.000 ;
    END
  END dyn0_dEo[55]
  PIN dyn0_dEo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END dyn0_dEo[56]
  PIN dyn0_dEo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 285.640 2500.000 286.240 ;
    END
  END dyn0_dEo[57]
  PIN dyn0_dEo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END dyn0_dEo[58]
  PIN dyn0_dEo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END dyn0_dEo[59]
  PIN dyn0_dEo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2216.840 2500.000 2217.440 ;
    END
  END dyn0_dEo[5]
  PIN dyn0_dEo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END dyn0_dEo[60]
  PIN dyn0_dEo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 2496.000 570.310 2500.000 ;
    END
  END dyn0_dEo[61]
  PIN dyn0_dEo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 2496.000 908.410 2500.000 ;
    END
  END dyn0_dEo[62]
  PIN dyn0_dEo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 693.640 2500.000 694.240 ;
    END
  END dyn0_dEo[63]
  PIN dyn0_dEo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2421.530 2496.000 2421.810 2500.000 ;
    END
  END dyn0_dEo[6]
  PIN dyn0_dEo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END dyn0_dEo[7]
  PIN dyn0_dEo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END dyn0_dEo[8]
  PIN dyn0_dEo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1985.640 4.000 1986.240 ;
    END
  END dyn0_dEo[9]
  PIN dyn0_dEo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.530 0.000 2260.810 4.000 ;
    END
  END dyn0_dEo_valid
  PIN dyn0_dEo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END dyn0_dEo_yummy
  PIN dyn0_dNo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.840 4.000 1469.440 ;
    END
  END dyn0_dNo[0]
  PIN dyn0_dNo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 2496.000 164.590 2500.000 ;
    END
  END dyn0_dNo[10]
  PIN dyn0_dNo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 2496.000 502.690 2500.000 ;
    END
  END dyn0_dNo[11]
  PIN dyn0_dNo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.450 0.000 2215.730 4.000 ;
    END
  END dyn0_dNo[12]
  PIN dyn0_dNo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.610 2496.000 2144.890 2500.000 ;
    END
  END dyn0_dNo[13]
  PIN dyn0_dNo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1829.240 2500.000 1829.840 ;
    END
  END dyn0_dNo[14]
  PIN dyn0_dNo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END dyn0_dNo[15]
  PIN dyn0_dNo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.890 2496.000 2383.170 2500.000 ;
    END
  END dyn0_dNo[16]
  PIN dyn0_dNo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2145.440 4.000 2146.040 ;
    END
  END dyn0_dNo[17]
  PIN dyn0_dNo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1404.240 2500.000 1404.840 ;
    END
  END dyn0_dNo[18]
  PIN dyn0_dNo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2349.440 4.000 2350.040 ;
    END
  END dyn0_dNo[19]
  PIN dyn0_dNo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 2496.000 1958.130 2500.000 ;
    END
  END dyn0_dNo[1]
  PIN dyn0_dNo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1040.440 2500.000 1041.040 ;
    END
  END dyn0_dNo[20]
  PIN dyn0_dNo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 2496.000 1159.570 2500.000 ;
    END
  END dyn0_dNo[21]
  PIN dyn0_dNo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 652.840 2500.000 653.440 ;
    END
  END dyn0_dNo[22]
  PIN dyn0_dNo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END dyn0_dNo[23]
  PIN dyn0_dNo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1655.840 2500.000 1656.440 ;
    END
  END dyn0_dNo[24]
  PIN dyn0_dNo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1873.440 2500.000 1874.040 ;
    END
  END dyn0_dNo[25]
  PIN dyn0_dNo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 2496.000 119.510 2500.000 ;
    END
  END dyn0_dNo[26]
  PIN dyn0_dNo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 0.000 1913.050 4.000 ;
    END
  END dyn0_dNo[27]
  PIN dyn0_dNo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2485.440 4.000 2486.040 ;
    END
  END dyn0_dNo[28]
  PIN dyn0_dNo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2050.240 2500.000 2050.840 ;
    END
  END dyn0_dNo[29]
  PIN dyn0_dNo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1193.440 2500.000 1194.040 ;
    END
  END dyn0_dNo[2]
  PIN dyn0_dNo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 0.000 2148.110 4.000 ;
    END
  END dyn0_dNo[30]
  PIN dyn0_dNo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2498.810 2496.000 2499.090 2500.000 ;
    END
  END dyn0_dNo[31]
  PIN dyn0_dNo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END dyn0_dNo[32]
  PIN dyn0_dNo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END dyn0_dNo[33]
  PIN dyn0_dNo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END dyn0_dNo[34]
  PIN dyn0_dNo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END dyn0_dNo[35]
  PIN dyn0_dNo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 598.440 2500.000 599.040 ;
    END
  END dyn0_dNo[36]
  PIN dyn0_dNo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 0.000 2103.030 4.000 ;
    END
  END dyn0_dNo[37]
  PIN dyn0_dNo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END dyn0_dNo[38]
  PIN dyn0_dNo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END dyn0_dNo[39]
  PIN dyn0_dNo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.890 2496.000 2222.170 2500.000 ;
    END
  END dyn0_dNo[3]
  PIN dyn0_dNo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 2496.000 1446.150 2500.000 ;
    END
  END dyn0_dNo[40]
  PIN dyn0_dNo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2199.840 2500.000 2200.440 ;
    END
  END dyn0_dNo[41]
  PIN dyn0_dNo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 2496.000 1645.790 2500.000 ;
    END
  END dyn0_dNo[42]
  PIN dyn0_dNo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 2496.000 1294.810 2500.000 ;
    END
  END dyn0_dNo[43]
  PIN dyn0_dNo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.650 2496.000 1925.930 2500.000 ;
    END
  END dyn0_dNo[44]
  PIN dyn0_dNo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END dyn0_dNo[45]
  PIN dyn0_dNo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 2496.000 2064.390 2500.000 ;
    END
  END dyn0_dNo[46]
  PIN dyn0_dNo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END dyn0_dNo[47]
  PIN dyn0_dNo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 2496.000 666.910 2500.000 ;
    END
  END dyn0_dNo[48]
  PIN dyn0_dNo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END dyn0_dNo[49]
  PIN dyn0_dNo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 4.000 ;
    END
  END dyn0_dNo[4]
  PIN dyn0_dNo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 292.440 2500.000 293.040 ;
    END
  END dyn0_dNo[50]
  PIN dyn0_dNo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 2496.000 232.210 2500.000 ;
    END
  END dyn0_dNo[51]
  PIN dyn0_dNo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END dyn0_dNo[52]
  PIN dyn0_dNo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END dyn0_dNo[53]
  PIN dyn0_dNo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2186.240 2500.000 2186.840 ;
    END
  END dyn0_dNo[54]
  PIN dyn0_dNo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 561.040 2500.000 561.640 ;
    END
  END dyn0_dNo[55]
  PIN dyn0_dNo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 2496.000 1983.890 2500.000 ;
    END
  END dyn0_dNo[56]
  PIN dyn0_dNo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END dyn0_dNo[57]
  PIN dyn0_dNo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1003.040 2500.000 1003.640 ;
    END
  END dyn0_dNo[58]
  PIN dyn0_dNo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 0.000 1848.650 4.000 ;
    END
  END dyn0_dNo[59]
  PIN dyn0_dNo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END dyn0_dNo[5]
  PIN dyn0_dNo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 2496.000 1120.930 2500.000 ;
    END
  END dyn0_dNo[60]
  PIN dyn0_dNo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.570 0.000 2363.850 4.000 ;
    END
  END dyn0_dNo[61]
  PIN dyn0_dNo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 0.000 2177.090 4.000 ;
    END
  END dyn0_dNo[62]
  PIN dyn0_dNo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 2496.000 1462.250 2500.000 ;
    END
  END dyn0_dNo[63]
  PIN dyn0_dNo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END dyn0_dNo[6]
  PIN dyn0_dNo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END dyn0_dNo[7]
  PIN dyn0_dNo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END dyn0_dNo[8]
  PIN dyn0_dNo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 2496.000 976.030 2500.000 ;
    END
  END dyn0_dNo[9]
  PIN dyn0_dNo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1842.840 2500.000 1843.440 ;
    END
  END dyn0_dNo_valid
  PIN dyn0_dNo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2498.810 0.000 2499.090 4.000 ;
    END
  END dyn0_dNo_yummy
  PIN dyn0_dSo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 2496.000 1655.450 2500.000 ;
    END
  END dyn0_dSo[0]
  PIN dyn0_dSo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1203.640 4.000 1204.240 ;
    END
  END dyn0_dSo[10]
  PIN dyn0_dSo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END dyn0_dSo[11]
  PIN dyn0_dSo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 2496.000 341.690 2500.000 ;
    END
  END dyn0_dSo[12]
  PIN dyn0_dSo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END dyn0_dSo[13]
  PIN dyn0_dSo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END dyn0_dSo[14]
  PIN dyn0_dSo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 2496.000 1555.630 2500.000 ;
    END
  END dyn0_dSo[15]
  PIN dyn0_dSo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.170 2496.000 1977.450 2500.000 ;
    END
  END dyn0_dSo[16]
  PIN dyn0_dSo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END dyn0_dSo[17]
  PIN dyn0_dSo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 2496.000 1175.670 2500.000 ;
    END
  END dyn0_dSo[18]
  PIN dyn0_dSo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 2496.000 1755.270 2500.000 ;
    END
  END dyn0_dSo[19]
  PIN dyn0_dSo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 958.840 2500.000 959.440 ;
    END
  END dyn0_dSo[1]
  PIN dyn0_dSo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 2496.000 541.330 2500.000 ;
    END
  END dyn0_dSo[20]
  PIN dyn0_dSo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1489.240 2500.000 1489.840 ;
    END
  END dyn0_dSo[21]
  PIN dyn0_dSo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 302.640 2500.000 303.240 ;
    END
  END dyn0_dSo[22]
  PIN dyn0_dSo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 2496.000 628.270 2500.000 ;
    END
  END dyn0_dSo[23]
  PIN dyn0_dSo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END dyn0_dSo[24]
  PIN dyn0_dSo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END dyn0_dSo[25]
  PIN dyn0_dSo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 778.640 2500.000 779.240 ;
    END
  END dyn0_dSo[26]
  PIN dyn0_dSo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 2496.000 1310.910 2500.000 ;
    END
  END dyn0_dSo[27]
  PIN dyn0_dSo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 2496.000 2312.330 2500.000 ;
    END
  END dyn0_dSo[28]
  PIN dyn0_dSo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END dyn0_dSo[29]
  PIN dyn0_dSo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.390 0.000 2302.670 4.000 ;
    END
  END dyn0_dSo[2]
  PIN dyn0_dSo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1016.640 2500.000 1017.240 ;
    END
  END dyn0_dSo[30]
  PIN dyn0_dSo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END dyn0_dSo[31]
  PIN dyn0_dSo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 2496.000 1375.310 2500.000 ;
    END
  END dyn0_dSo[32]
  PIN dyn0_dSo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1700.040 4.000 1700.640 ;
    END
  END dyn0_dSo[33]
  PIN dyn0_dSo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END dyn0_dSo[34]
  PIN dyn0_dSo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END dyn0_dSo[35]
  PIN dyn0_dSo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1356.640 2500.000 1357.240 ;
    END
  END dyn0_dSo[36]
  PIN dyn0_dSo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END dyn0_dSo[37]
  PIN dyn0_dSo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 2496.000 1027.550 2500.000 ;
    END
  END dyn0_dSo[38]
  PIN dyn0_dSo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END dyn0_dSo[39]
  PIN dyn0_dSo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END dyn0_dSo[3]
  PIN dyn0_dSo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END dyn0_dSo[40]
  PIN dyn0_dSo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1938.040 2500.000 1938.640 ;
    END
  END dyn0_dSo[41]
  PIN dyn0_dSo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.450 2496.000 2215.730 2500.000 ;
    END
  END dyn0_dSo[42]
  PIN dyn0_dSo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 2496.000 818.250 2500.000 ;
    END
  END dyn0_dSo[43]
  PIN dyn0_dSo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END dyn0_dSo[44]
  PIN dyn0_dSo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.150 2496.000 2167.430 2500.000 ;
    END
  END dyn0_dSo[45]
  PIN dyn0_dSo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 2496.000 1594.270 2500.000 ;
    END
  END dyn0_dSo[46]
  PIN dyn0_dSo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.990 2496.000 2238.270 2500.000 ;
    END
  END dyn0_dSo[47]
  PIN dyn0_dSo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END dyn0_dSo[48]
  PIN dyn0_dSo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 476.040 2500.000 476.640 ;
    END
  END dyn0_dSo[49]
  PIN dyn0_dSo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1346.440 2500.000 1347.040 ;
    END
  END dyn0_dSo[4]
  PIN dyn0_dSo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 2496.000 61.550 2500.000 ;
    END
  END dyn0_dSo[50]
  PIN dyn0_dSo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 2496.000 412.530 2500.000 ;
    END
  END dyn0_dSo[51]
  PIN dyn0_dSo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.450 2496.000 2054.730 2500.000 ;
    END
  END dyn0_dSo[52]
  PIN dyn0_dSo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 4.000 ;
    END
  END dyn0_dSo[53]
  PIN dyn0_dSo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 0.000 1272.270 4.000 ;
    END
  END dyn0_dSo[54]
  PIN dyn0_dSo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1798.640 2500.000 1799.240 ;
    END
  END dyn0_dSo[55]
  PIN dyn0_dSo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 265.240 2500.000 265.840 ;
    END
  END dyn0_dSo[56]
  PIN dyn0_dSo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2278.040 4.000 2278.640 ;
    END
  END dyn0_dSo[57]
  PIN dyn0_dSo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END dyn0_dSo[58]
  PIN dyn0_dSo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END dyn0_dSo[59]
  PIN dyn0_dSo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1159.440 2500.000 1160.040 ;
    END
  END dyn0_dSo[5]
  PIN dyn0_dSo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.590 0.000 2334.870 4.000 ;
    END
  END dyn0_dSo[60]
  PIN dyn0_dSo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 2496.000 1365.650 2500.000 ;
    END
  END dyn0_dSo[61]
  PIN dyn0_dSo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 2496.000 1523.430 2500.000 ;
    END
  END dyn0_dSo[62]
  PIN dyn0_dSo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 0.000 1220.750 4.000 ;
    END
  END dyn0_dSo[63]
  PIN dyn0_dSo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1659.240 2500.000 1659.840 ;
    END
  END dyn0_dSo[6]
  PIN dyn0_dSo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1788.440 2500.000 1789.040 ;
    END
  END dyn0_dSo[7]
  PIN dyn0_dSo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.510 0.000 1967.790 4.000 ;
    END
  END dyn0_dSo[8]
  PIN dyn0_dSo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END dyn0_dSo[9]
  PIN dyn0_dSo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2373.240 4.000 2373.840 ;
    END
  END dyn0_dSo_valid
  PIN dyn0_dSo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.670 2496.000 1896.950 2500.000 ;
    END
  END dyn0_dSo_yummy
  PIN dyn0_dWo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 278.840 2500.000 279.440 ;
    END
  END dyn0_dWo[0]
  PIN dyn0_dWo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.270 2496.000 2476.550 2500.000 ;
    END
  END dyn0_dWo[10]
  PIN dyn0_dWo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END dyn0_dWo[11]
  PIN dyn0_dWo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.510 2496.000 2128.790 2500.000 ;
    END
  END dyn0_dWo[12]
  PIN dyn0_dWo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 2496.000 1745.610 2500.000 ;
    END
  END dyn0_dWo[13]
  PIN dyn0_dWo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END dyn0_dWo[14]
  PIN dyn0_dWo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END dyn0_dWo[15]
  PIN dyn0_dWo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END dyn0_dWo[16]
  PIN dyn0_dWo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 924.840 2500.000 925.440 ;
    END
  END dyn0_dWo[17]
  PIN dyn0_dWo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 0.000 1133.810 4.000 ;
    END
  END dyn0_dWo[18]
  PIN dyn0_dWo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END dyn0_dWo[19]
  PIN dyn0_dWo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END dyn0_dWo[1]
  PIN dyn0_dWo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 2496.000 1098.390 2500.000 ;
    END
  END dyn0_dWo[20]
  PIN dyn0_dWo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2359.640 2500.000 2360.240 ;
    END
  END dyn0_dWo[21]
  PIN dyn0_dWo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 2496.000 2109.470 2500.000 ;
    END
  END dyn0_dWo[22]
  PIN dyn0_dWo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 2496.000 740.970 2500.000 ;
    END
  END dyn0_dWo[23]
  PIN dyn0_dWo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1421.240 2500.000 1421.840 ;
    END
  END dyn0_dWo[24]
  PIN dyn0_dWo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2403.840 4.000 2404.440 ;
    END
  END dyn0_dWo[25]
  PIN dyn0_dWo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.230 2496.000 2051.510 2500.000 ;
    END
  END dyn0_dWo[26]
  PIN dyn0_dWo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 2496.000 2212.510 2500.000 ;
    END
  END dyn0_dWo[27]
  PIN dyn0_dWo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 2496.000 344.910 2500.000 ;
    END
  END dyn0_dWo[28]
  PIN dyn0_dWo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2418.310 2496.000 2418.590 2500.000 ;
    END
  END dyn0_dWo[29]
  PIN dyn0_dWo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 2496.000 773.170 2500.000 ;
    END
  END dyn0_dWo[2]
  PIN dyn0_dWo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END dyn0_dWo[30]
  PIN dyn0_dWo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2369.840 4.000 2370.440 ;
    END
  END dyn0_dWo[31]
  PIN dyn0_dWo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 88.440 2500.000 89.040 ;
    END
  END dyn0_dWo[32]
  PIN dyn0_dWo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END dyn0_dWo[33]
  PIN dyn0_dWo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END dyn0_dWo[34]
  PIN dyn0_dWo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1948.240 2500.000 1948.840 ;
    END
  END dyn0_dWo[35]
  PIN dyn0_dWo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.040 4.000 1394.640 ;
    END
  END dyn0_dWo[36]
  PIN dyn0_dWo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 707.240 2500.000 707.840 ;
    END
  END dyn0_dWo[37]
  PIN dyn0_dWo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END dyn0_dWo[38]
  PIN dyn0_dWo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END dyn0_dWo[39]
  PIN dyn0_dWo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1785.040 2500.000 1785.640 ;
    END
  END dyn0_dWo[3]
  PIN dyn0_dWo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 2496.000 1607.150 2500.000 ;
    END
  END dyn0_dWo[40]
  PIN dyn0_dWo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END dyn0_dWo[41]
  PIN dyn0_dWo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END dyn0_dWo[42]
  PIN dyn0_dWo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1876.840 2500.000 1877.440 ;
    END
  END dyn0_dWo[43]
  PIN dyn0_dWo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 0.000 1874.410 4.000 ;
    END
  END dyn0_dWo[44]
  PIN dyn0_dWo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 4.000 ;
    END
  END dyn0_dWo[45]
  PIN dyn0_dWo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2380.040 2500.000 2380.640 ;
    END
  END dyn0_dWo[46]
  PIN dyn0_dWo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END dyn0_dWo[47]
  PIN dyn0_dWo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END dyn0_dWo[48]
  PIN dyn0_dWo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1795.240 4.000 1795.840 ;
    END
  END dyn0_dWo[49]
  PIN dyn0_dWo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1931.240 2500.000 1931.840 ;
    END
  END dyn0_dWo[4]
  PIN dyn0_dWo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 2496.000 930.950 2500.000 ;
    END
  END dyn0_dWo[50]
  PIN dyn0_dWo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END dyn0_dWo[51]
  PIN dyn0_dWo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 2496.000 286.950 2500.000 ;
    END
  END dyn0_dWo[52]
  PIN dyn0_dWo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 2496.000 45.450 2500.000 ;
    END
  END dyn0_dWo[53]
  PIN dyn0_dWo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1859.840 2500.000 1860.440 ;
    END
  END dyn0_dWo[54]
  PIN dyn0_dWo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2087.640 2500.000 2088.240 ;
    END
  END dyn0_dWo[55]
  PIN dyn0_dWo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 2496.000 647.590 2500.000 ;
    END
  END dyn0_dWo[56]
  PIN dyn0_dWo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END dyn0_dWo[57]
  PIN dyn0_dWo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.810 2496.000 2338.090 2500.000 ;
    END
  END dyn0_dWo[58]
  PIN dyn0_dWo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END dyn0_dWo[59]
  PIN dyn0_dWo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END dyn0_dWo[5]
  PIN dyn0_dWo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END dyn0_dWo[60]
  PIN dyn0_dWo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 2496.000 2392.830 2500.000 ;
    END
  END dyn0_dWo[61]
  PIN dyn0_dWo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2128.440 4.000 2129.040 ;
    END
  END dyn0_dWo[62]
  PIN dyn0_dWo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 2496.000 299.830 2500.000 ;
    END
  END dyn0_dWo[63]
  PIN dyn0_dWo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1241.040 2500.000 1241.640 ;
    END
  END dyn0_dWo[6]
  PIN dyn0_dWo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 367.240 2500.000 367.840 ;
    END
  END dyn0_dWo[7]
  PIN dyn0_dWo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END dyn0_dWo[8]
  PIN dyn0_dWo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END dyn0_dWo[9]
  PIN dyn0_dWo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END dyn0_dWo_valid
  PIN dyn0_dWo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1771.440 2500.000 1772.040 ;
    END
  END dyn0_dWo_yummy
  PIN dyn0_dataIn_E[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END dyn0_dataIn_E[0]
  PIN dyn0_dataIn_E[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 0.000 1723.070 4.000 ;
    END
  END dyn0_dataIn_E[10]
  PIN dyn0_dataIn_E[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 0.000 1900.170 4.000 ;
    END
  END dyn0_dataIn_E[11]
  PIN dyn0_dataIn_E[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END dyn0_dataIn_E[12]
  PIN dyn0_dataIn_E[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 0.000 2115.910 4.000 ;
    END
  END dyn0_dataIn_E[13]
  PIN dyn0_dataIn_E[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 584.840 2500.000 585.440 ;
    END
  END dyn0_dataIn_E[14]
  PIN dyn0_dataIn_E[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 2496.000 151.710 2500.000 ;
    END
  END dyn0_dataIn_E[15]
  PIN dyn0_dataIn_E[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 2496.000 1574.950 2500.000 ;
    END
  END dyn0_dataIn_E[16]
  PIN dyn0_dataIn_E[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END dyn0_dataIn_E[17]
  PIN dyn0_dataIn_E[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END dyn0_dataIn_E[18]
  PIN dyn0_dataIn_E[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.670 0.000 2379.950 4.000 ;
    END
  END dyn0_dataIn_E[19]
  PIN dyn0_dataIn_E[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 2496.000 779.610 2500.000 ;
    END
  END dyn0_dataIn_E[1]
  PIN dyn0_dataIn_E[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END dyn0_dataIn_E[20]
  PIN dyn0_dataIn_E[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END dyn0_dataIn_E[21]
  PIN dyn0_dataIn_E[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END dyn0_dataIn_E[22]
  PIN dyn0_dataIn_E[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 200.640 2500.000 201.240 ;
    END
  END dyn0_dataIn_E[23]
  PIN dyn0_dataIn_E[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 2496.000 1558.850 2500.000 ;
    END
  END dyn0_dataIn_E[24]
  PIN dyn0_dataIn_E[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 2496.000 19.690 2500.000 ;
    END
  END dyn0_dataIn_E[25]
  PIN dyn0_dataIn_E[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 20.440 2500.000 21.040 ;
    END
  END dyn0_dataIn_E[26]
  PIN dyn0_dataIn_E[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 0.000 2109.470 4.000 ;
    END
  END dyn0_dataIn_E[27]
  PIN dyn0_dataIn_E[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END dyn0_dataIn_E[28]
  PIN dyn0_dataIn_E[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1771.440 4.000 1772.040 ;
    END
  END dyn0_dataIn_E[29]
  PIN dyn0_dataIn_E[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END dyn0_dataIn_E[2]
  PIN dyn0_dataIn_E[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1288.640 2500.000 1289.240 ;
    END
  END dyn0_dataIn_E[30]
  PIN dyn0_dataIn_E[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1441.640 2500.000 1442.240 ;
    END
  END dyn0_dataIn_E[31]
  PIN dyn0_dataIn_E[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 2496.000 1085.510 2500.000 ;
    END
  END dyn0_dataIn_E[32]
  PIN dyn0_dataIn_E[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2346.040 4.000 2346.640 ;
    END
  END dyn0_dataIn_E[33]
  PIN dyn0_dataIn_E[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.870 2496.000 2251.150 2500.000 ;
    END
  END dyn0_dataIn_E[34]
  PIN dyn0_dataIn_E[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END dyn0_dataIn_E[35]
  PIN dyn0_dataIn_E[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END dyn0_dataIn_E[36]
  PIN dyn0_dataIn_E[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 2496.000 673.350 2500.000 ;
    END
  END dyn0_dataIn_E[37]
  PIN dyn0_dataIn_E[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1975.440 4.000 1976.040 ;
    END
  END dyn0_dataIn_E[38]
  PIN dyn0_dataIn_E[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END dyn0_dataIn_E[39]
  PIN dyn0_dataIn_E[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 2496.000 100.190 2500.000 ;
    END
  END dyn0_dataIn_E[3]
  PIN dyn0_dataIn_E[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END dyn0_dataIn_E[40]
  PIN dyn0_dataIn_E[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 2496.000 1900.170 2500.000 ;
    END
  END dyn0_dataIn_E[41]
  PIN dyn0_dataIn_E[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.710 0.000 2321.990 4.000 ;
    END
  END dyn0_dataIn_E[42]
  PIN dyn0_dataIn_E[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.830 0.000 2309.110 4.000 ;
    END
  END dyn0_dataIn_E[43]
  PIN dyn0_dataIn_E[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END dyn0_dataIn_E[44]
  PIN dyn0_dataIn_E[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END dyn0_dataIn_E[45]
  PIN dyn0_dataIn_E[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 0.000 1880.850 4.000 ;
    END
  END dyn0_dataIn_E[46]
  PIN dyn0_dataIn_E[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 2496.000 966.370 2500.000 ;
    END
  END dyn0_dataIn_E[47]
  PIN dyn0_dataIn_E[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 856.840 2500.000 857.440 ;
    END
  END dyn0_dataIn_E[48]
  PIN dyn0_dataIn_E[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 846.640 2500.000 847.240 ;
    END
  END dyn0_dataIn_E[49]
  PIN dyn0_dataIn_E[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1570.840 4.000 1571.440 ;
    END
  END dyn0_dataIn_E[4]
  PIN dyn0_dataIn_E[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END dyn0_dataIn_E[50]
  PIN dyn0_dataIn_E[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2461.640 2500.000 2462.240 ;
    END
  END dyn0_dataIn_E[51]
  PIN dyn0_dataIn_E[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 2496.000 132.390 2500.000 ;
    END
  END dyn0_dataIn_E[52]
  PIN dyn0_dataIn_E[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1642.240 4.000 1642.840 ;
    END
  END dyn0_dataIn_E[53]
  PIN dyn0_dataIn_E[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 2496.000 135.610 2500.000 ;
    END
  END dyn0_dataIn_E[54]
  PIN dyn0_dataIn_E[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1088.040 2500.000 1088.640 ;
    END
  END dyn0_dataIn_E[55]
  PIN dyn0_dataIn_E[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 2496.000 927.730 2500.000 ;
    END
  END dyn0_dataIn_E[56]
  PIN dyn0_dataIn_E[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 319.640 2500.000 320.240 ;
    END
  END dyn0_dataIn_E[57]
  PIN dyn0_dataIn_E[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2131.840 4.000 2132.440 ;
    END
  END dyn0_dataIn_E[58]
  PIN dyn0_dataIn_E[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 744.640 2500.000 745.240 ;
    END
  END dyn0_dataIn_E[59]
  PIN dyn0_dataIn_E[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END dyn0_dataIn_E[5]
  PIN dyn0_dataIn_E[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 853.440 2500.000 854.040 ;
    END
  END dyn0_dataIn_E[60]
  PIN dyn0_dataIn_E[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.840 4.000 1316.440 ;
    END
  END dyn0_dataIn_E[61]
  PIN dyn0_dataIn_E[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1564.040 2500.000 1564.640 ;
    END
  END dyn0_dataIn_E[62]
  PIN dyn0_dataIn_E[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END dyn0_dataIn_E[63]
  PIN dyn0_dataIn_E[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1897.240 2500.000 1897.840 ;
    END
  END dyn0_dataIn_E[6]
  PIN dyn0_dataIn_E[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2074.040 2500.000 2074.640 ;
    END
  END dyn0_dataIn_E[7]
  PIN dyn0_dataIn_E[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END dyn0_dataIn_E[8]
  PIN dyn0_dataIn_E[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 176.840 2500.000 177.440 ;
    END
  END dyn0_dataIn_E[9]
  PIN dyn0_dataIn_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 2496.000 409.310 2500.000 ;
    END
  END dyn0_dataIn_N[0]
  PIN dyn0_dataIn_N[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 2496.000 203.230 2500.000 ;
    END
  END dyn0_dataIn_N[10]
  PIN dyn0_dataIn_N[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1812.240 2500.000 1812.840 ;
    END
  END dyn0_dataIn_N[11]
  PIN dyn0_dataIn_N[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 0.000 1591.050 4.000 ;
    END
  END dyn0_dataIn_N[12]
  PIN dyn0_dataIn_N[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2454.840 2500.000 2455.440 ;
    END
  END dyn0_dataIn_N[13]
  PIN dyn0_dataIn_N[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 646.040 2500.000 646.640 ;
    END
  END dyn0_dataIn_N[14]
  PIN dyn0_dataIn_N[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 2496.000 103.410 2500.000 ;
    END
  END dyn0_dataIn_N[15]
  PIN dyn0_dataIn_N[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END dyn0_dataIn_N[16]
  PIN dyn0_dataIn_N[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END dyn0_dataIn_N[17]
  PIN dyn0_dataIn_N[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 2496.000 1178.890 2500.000 ;
    END
  END dyn0_dataIn_N[18]
  PIN dyn0_dataIn_N[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1332.840 2500.000 1333.440 ;
    END
  END dyn0_dataIn_N[19]
  PIN dyn0_dataIn_N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END dyn0_dataIn_N[1]
  PIN dyn0_dataIn_N[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END dyn0_dataIn_N[20]
  PIN dyn0_dataIn_N[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 2496.000 731.310 2500.000 ;
    END
  END dyn0_dataIn_N[21]
  PIN dyn0_dataIn_N[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2264.440 2500.000 2265.040 ;
    END
  END dyn0_dataIn_N[22]
  PIN dyn0_dataIn_N[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END dyn0_dataIn_N[23]
  PIN dyn0_dataIn_N[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 0.000 1706.970 4.000 ;
    END
  END dyn0_dataIn_N[24]
  PIN dyn0_dataIn_N[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 2496.000 1391.410 2500.000 ;
    END
  END dyn0_dataIn_N[25]
  PIN dyn0_dataIn_N[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1853.040 2500.000 1853.640 ;
    END
  END dyn0_dataIn_N[26]
  PIN dyn0_dataIn_N[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1349.840 2500.000 1350.440 ;
    END
  END dyn0_dataIn_N[27]
  PIN dyn0_dataIn_N[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END dyn0_dataIn_N[28]
  PIN dyn0_dataIn_N[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2359.640 4.000 2360.240 ;
    END
  END dyn0_dataIn_N[29]
  PIN dyn0_dataIn_N[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END dyn0_dataIn_N[2]
  PIN dyn0_dataIn_N[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END dyn0_dataIn_N[30]
  PIN dyn0_dataIn_N[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 2496.000 1204.650 2500.000 ;
    END
  END dyn0_dataIn_N[31]
  PIN dyn0_dataIn_N[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 2496.000 1156.350 2500.000 ;
    END
  END dyn0_dataIn_N[32]
  PIN dyn0_dataIn_N[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 482.840 2500.000 483.440 ;
    END
  END dyn0_dataIn_N[33]
  PIN dyn0_dataIn_N[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2084.240 4.000 2084.840 ;
    END
  END dyn0_dataIn_N[34]
  PIN dyn0_dataIn_N[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 2496.000 383.550 2500.000 ;
    END
  END dyn0_dataIn_N[35]
  PIN dyn0_dataIn_N[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1326.040 2500.000 1326.640 ;
    END
  END dyn0_dataIn_N[36]
  PIN dyn0_dataIn_N[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 2496.000 1127.370 2500.000 ;
    END
  END dyn0_dataIn_N[37]
  PIN dyn0_dataIn_N[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 2496.000 309.490 2500.000 ;
    END
  END dyn0_dataIn_N[38]
  PIN dyn0_dataIn_N[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 469.240 2500.000 469.840 ;
    END
  END dyn0_dataIn_N[39]
  PIN dyn0_dataIn_N[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 2496.000 2080.490 2500.000 ;
    END
  END dyn0_dataIn_N[3]
  PIN dyn0_dataIn_N[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.470 2496.000 2025.750 2500.000 ;
    END
  END dyn0_dataIn_N[40]
  PIN dyn0_dataIn_N[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 465.840 2500.000 466.440 ;
    END
  END dyn0_dataIn_N[41]
  PIN dyn0_dataIn_N[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.730 2496.000 2132.010 2500.000 ;
    END
  END dyn0_dataIn_N[42]
  PIN dyn0_dataIn_N[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END dyn0_dataIn_N[43]
  PIN dyn0_dataIn_N[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 2496.000 1275.490 2500.000 ;
    END
  END dyn0_dataIn_N[44]
  PIN dyn0_dataIn_N[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1468.840 2500.000 1469.440 ;
    END
  END dyn0_dataIn_N[45]
  PIN dyn0_dataIn_N[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2308.640 4.000 2309.240 ;
    END
  END dyn0_dataIn_N[46]
  PIN dyn0_dataIn_N[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2400.440 4.000 2401.040 ;
    END
  END dyn0_dataIn_N[47]
  PIN dyn0_dataIn_N[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 2496.000 364.230 2500.000 ;
    END
  END dyn0_dataIn_N[48]
  PIN dyn0_dataIn_N[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 2496.000 303.050 2500.000 ;
    END
  END dyn0_dataIn_N[49]
  PIN dyn0_dataIn_N[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 816.040 2500.000 816.640 ;
    END
  END dyn0_dataIn_N[4]
  PIN dyn0_dataIn_N[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 241.440 2500.000 242.040 ;
    END
  END dyn0_dataIn_N[50]
  PIN dyn0_dataIn_N[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1615.040 2500.000 1615.640 ;
    END
  END dyn0_dataIn_N[51]
  PIN dyn0_dataIn_N[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1550.440 2500.000 1551.040 ;
    END
  END dyn0_dataIn_N[52]
  PIN dyn0_dataIn_N[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END dyn0_dataIn_N[53]
  PIN dyn0_dataIn_N[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.840 4.000 1673.440 ;
    END
  END dyn0_dataIn_N[54]
  PIN dyn0_dataIn_N[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END dyn0_dataIn_N[55]
  PIN dyn0_dataIn_N[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END dyn0_dataIn_N[56]
  PIN dyn0_dataIn_N[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1958.440 4.000 1959.040 ;
    END
  END dyn0_dataIn_N[57]
  PIN dyn0_dataIn_N[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1628.640 2500.000 1629.240 ;
    END
  END dyn0_dataIn_N[58]
  PIN dyn0_dataIn_N[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1914.240 2500.000 1914.840 ;
    END
  END dyn0_dataIn_N[59]
  PIN dyn0_dataIn_N[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 720.840 2500.000 721.440 ;
    END
  END dyn0_dataIn_N[5]
  PIN dyn0_dataIn_N[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 982.640 2500.000 983.240 ;
    END
  END dyn0_dataIn_N[60]
  PIN dyn0_dataIn_N[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 323.040 2500.000 323.640 ;
    END
  END dyn0_dataIn_N[61]
  PIN dyn0_dataIn_N[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END dyn0_dataIn_N[62]
  PIN dyn0_dataIn_N[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1547.040 2500.000 1547.640 ;
    END
  END dyn0_dataIn_N[63]
  PIN dyn0_dataIn_N[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1717.040 2500.000 1717.640 ;
    END
  END dyn0_dataIn_N[6]
  PIN dyn0_dataIn_N[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 2496.000 953.490 2500.000 ;
    END
  END dyn0_dataIn_N[7]
  PIN dyn0_dataIn_N[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2108.040 2500.000 2108.640 ;
    END
  END dyn0_dataIn_N[8]
  PIN dyn0_dataIn_N[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END dyn0_dataIn_N[9]
  PIN dyn0_dataIn_S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END dyn0_dataIn_S[0]
  PIN dyn0_dataIn_S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2257.640 4.000 2258.240 ;
    END
  END dyn0_dataIn_S[10]
  PIN dyn0_dataIn_S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 588.240 2500.000 588.840 ;
    END
  END dyn0_dataIn_S[11]
  PIN dyn0_dataIn_S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 2496.000 464.050 2500.000 ;
    END
  END dyn0_dataIn_S[12]
  PIN dyn0_dataIn_S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END dyn0_dataIn_S[13]
  PIN dyn0_dataIn_S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.410 0.000 2273.690 4.000 ;
    END
  END dyn0_dataIn_S[14]
  PIN dyn0_dataIn_S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2291.640 4.000 2292.240 ;
    END
  END dyn0_dataIn_S[15]
  PIN dyn0_dataIn_S[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 0.000 1610.370 4.000 ;
    END
  END dyn0_dataIn_S[16]
  PIN dyn0_dataIn_S[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.710 2496.000 1999.990 2500.000 ;
    END
  END dyn0_dataIn_S[17]
  PIN dyn0_dataIn_S[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 578.040 2500.000 578.640 ;
    END
  END dyn0_dataIn_S[18]
  PIN dyn0_dataIn_S[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 0.000 1710.190 4.000 ;
    END
  END dyn0_dataIn_S[19]
  PIN dyn0_dataIn_S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END dyn0_dataIn_S[1]
  PIN dyn0_dataIn_S[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2114.840 2500.000 2115.440 ;
    END
  END dyn0_dataIn_S[20]
  PIN dyn0_dataIn_S[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2267.840 4.000 2268.440 ;
    END
  END dyn0_dataIn_S[21]
  PIN dyn0_dataIn_S[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 0.000 2086.930 4.000 ;
    END
  END dyn0_dataIn_S[22]
  PIN dyn0_dataIn_S[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 2496.000 1249.730 2500.000 ;
    END
  END dyn0_dataIn_S[23]
  PIN dyn0_dataIn_S[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 2496.000 158.150 2500.000 ;
    END
  END dyn0_dataIn_S[24]
  PIN dyn0_dataIn_S[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 2496.000 1459.030 2500.000 ;
    END
  END dyn0_dataIn_S[25]
  PIN dyn0_dataIn_S[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END dyn0_dataIn_S[26]
  PIN dyn0_dataIn_S[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 829.640 2500.000 830.240 ;
    END
  END dyn0_dataIn_S[27]
  PIN dyn0_dataIn_S[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END dyn0_dataIn_S[28]
  PIN dyn0_dataIn_S[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.770 2496.000 2235.050 2500.000 ;
    END
  END dyn0_dataIn_S[29]
  PIN dyn0_dataIn_S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END dyn0_dataIn_S[2]
  PIN dyn0_dataIn_S[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 2496.000 734.530 2500.000 ;
    END
  END dyn0_dataIn_S[30]
  PIN dyn0_dataIn_S[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 2496.000 87.310 2500.000 ;
    END
  END dyn0_dataIn_S[31]
  PIN dyn0_dataIn_S[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 2496.000 1072.630 2500.000 ;
    END
  END dyn0_dataIn_S[32]
  PIN dyn0_dataIn_S[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1043.840 2500.000 1044.440 ;
    END
  END dyn0_dataIn_S[33]
  PIN dyn0_dataIn_S[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END dyn0_dataIn_S[34]
  PIN dyn0_dataIn_S[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END dyn0_dataIn_S[35]
  PIN dyn0_dataIn_S[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END dyn0_dataIn_S[36]
  PIN dyn0_dataIn_S[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END dyn0_dataIn_S[37]
  PIN dyn0_dataIn_S[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 2496.000 721.650 2500.000 ;
    END
  END dyn0_dataIn_S[38]
  PIN dyn0_dataIn_S[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 2496.000 1149.910 2500.000 ;
    END
  END dyn0_dataIn_S[39]
  PIN dyn0_dataIn_S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1839.440 2500.000 1840.040 ;
    END
  END dyn0_dataIn_S[3]
  PIN dyn0_dataIn_S[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1890.440 4.000 1891.040 ;
    END
  END dyn0_dataIn_S[40]
  PIN dyn0_dataIn_S[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 0.000 2212.510 4.000 ;
    END
  END dyn0_dataIn_S[41]
  PIN dyn0_dataIn_S[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 2496.000 934.170 2500.000 ;
    END
  END dyn0_dataIn_S[42]
  PIN dyn0_dataIn_S[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 775.240 2500.000 775.840 ;
    END
  END dyn0_dataIn_S[43]
  PIN dyn0_dataIn_S[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 2496.000 2122.350 2500.000 ;
    END
  END dyn0_dataIn_S[44]
  PIN dyn0_dataIn_S[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.970 0.000 2267.250 4.000 ;
    END
  END dyn0_dataIn_S[45]
  PIN dyn0_dataIn_S[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END dyn0_dataIn_S[46]
  PIN dyn0_dataIn_S[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1594.640 2500.000 1595.240 ;
    END
  END dyn0_dataIn_S[47]
  PIN dyn0_dataIn_S[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.150 0.000 2006.430 4.000 ;
    END
  END dyn0_dataIn_S[48]
  PIN dyn0_dataIn_S[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.840 4.000 1758.440 ;
    END
  END dyn0_dataIn_S[49]
  PIN dyn0_dataIn_S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END dyn0_dataIn_S[4]
  PIN dyn0_dataIn_S[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2427.640 2500.000 2428.240 ;
    END
  END dyn0_dataIn_S[50]
  PIN dyn0_dataIn_S[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END dyn0_dataIn_S[51]
  PIN dyn0_dataIn_S[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 2496.000 2396.050 2500.000 ;
    END
  END dyn0_dataIn_S[52]
  PIN dyn0_dataIn_S[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2233.840 4.000 2234.440 ;
    END
  END dyn0_dataIn_S[53]
  PIN dyn0_dataIn_S[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 255.040 2500.000 255.640 ;
    END
  END dyn0_dataIn_S[54]
  PIN dyn0_dataIn_S[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 690.240 2500.000 690.840 ;
    END
  END dyn0_dataIn_S[55]
  PIN dyn0_dataIn_S[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END dyn0_dataIn_S[56]
  PIN dyn0_dataIn_S[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.270 0.000 1993.550 4.000 ;
    END
  END dyn0_dataIn_S[57]
  PIN dyn0_dataIn_S[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2261.040 4.000 2261.640 ;
    END
  END dyn0_dataIn_S[58]
  PIN dyn0_dataIn_S[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END dyn0_dataIn_S[59]
  PIN dyn0_dataIn_S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 952.040 2500.000 952.640 ;
    END
  END dyn0_dataIn_S[5]
  PIN dyn0_dataIn_S[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END dyn0_dataIn_S[60]
  PIN dyn0_dataIn_S[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1553.840 2500.000 1554.440 ;
    END
  END dyn0_dataIn_S[61]
  PIN dyn0_dataIn_S[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 0.000 1301.250 4.000 ;
    END
  END dyn0_dataIn_S[62]
  PIN dyn0_dataIn_S[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1710.240 2500.000 1710.840 ;
    END
  END dyn0_dataIn_S[63]
  PIN dyn0_dataIn_S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END dyn0_dataIn_S[6]
  PIN dyn0_dataIn_S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 2496.000 167.810 2500.000 ;
    END
  END dyn0_dataIn_S[7]
  PIN dyn0_dataIn_S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 2496.000 1539.530 2500.000 ;
    END
  END dyn0_dataIn_S[8]
  PIN dyn0_dataIn_S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2189.640 4.000 2190.240 ;
    END
  END dyn0_dataIn_S[9]
  PIN dyn0_dataIn_W[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.190 0.000 1626.470 4.000 ;
    END
  END dyn0_dataIn_W[0]
  PIN dyn0_dataIn_W[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 2496.000 2106.250 2500.000 ;
    END
  END dyn0_dataIn_W[10]
  PIN dyn0_dataIn_W[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END dyn0_dataIn_W[11]
  PIN dyn0_dataIn_W[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.690 2496.000 2028.970 2500.000 ;
    END
  END dyn0_dataIn_W[12]
  PIN dyn0_dataIn_W[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 2496.000 154.930 2500.000 ;
    END
  END dyn0_dataIn_W[13]
  PIN dyn0_dataIn_W[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 2496.000 1536.310 2500.000 ;
    END
  END dyn0_dataIn_W[14]
  PIN dyn0_dataIn_W[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 2496.000 1223.970 2500.000 ;
    END
  END dyn0_dataIn_W[15]
  PIN dyn0_dataIn_W[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END dyn0_dataIn_W[16]
  PIN dyn0_dataIn_W[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 2496.000 1758.490 2500.000 ;
    END
  END dyn0_dataIn_W[17]
  PIN dyn0_dataIn_W[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1999.240 2500.000 1999.840 ;
    END
  END dyn0_dataIn_W[18]
  PIN dyn0_dataIn_W[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 2496.000 1890.510 2500.000 ;
    END
  END dyn0_dataIn_W[19]
  PIN dyn0_dataIn_W[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 2496.000 1652.230 2500.000 ;
    END
  END dyn0_dataIn_W[1]
  PIN dyn0_dataIn_W[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 37.440 2500.000 38.040 ;
    END
  END dyn0_dataIn_W[20]
  PIN dyn0_dataIn_W[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2427.640 4.000 2428.240 ;
    END
  END dyn0_dataIn_W[21]
  PIN dyn0_dataIn_W[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 275.440 2500.000 276.040 ;
    END
  END dyn0_dataIn_W[22]
  PIN dyn0_dataIn_W[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 0.000 2396.050 4.000 ;
    END
  END dyn0_dataIn_W[23]
  PIN dyn0_dataIn_W[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.450 2496.000 2376.730 2500.000 ;
    END
  END dyn0_dataIn_W[24]
  PIN dyn0_dataIn_W[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 2496.000 1706.970 2500.000 ;
    END
  END dyn0_dataIn_W[25]
  PIN dyn0_dataIn_W[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 2496.000 985.690 2500.000 ;
    END
  END dyn0_dataIn_W[26]
  PIN dyn0_dataIn_W[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1703.440 4.000 1704.040 ;
    END
  END dyn0_dataIn_W[27]
  PIN dyn0_dataIn_W[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2271.240 2500.000 2271.840 ;
    END
  END dyn0_dataIn_W[28]
  PIN dyn0_dataIn_W[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.510 0.000 2289.790 4.000 ;
    END
  END dyn0_dataIn_W[29]
  PIN dyn0_dataIn_W[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1424.640 2500.000 1425.240 ;
    END
  END dyn0_dataIn_W[2]
  PIN dyn0_dataIn_W[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1224.040 2500.000 1224.640 ;
    END
  END dyn0_dataIn_W[30]
  PIN dyn0_dataIn_W[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END dyn0_dataIn_W[31]
  PIN dyn0_dataIn_W[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.370 0.000 2492.650 4.000 ;
    END
  END dyn0_dataIn_W[32]
  PIN dyn0_dataIn_W[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1618.440 4.000 1619.040 ;
    END
  END dyn0_dataIn_W[33]
  PIN dyn0_dataIn_W[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 0.000 1549.190 4.000 ;
    END
  END dyn0_dataIn_W[34]
  PIN dyn0_dataIn_W[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END dyn0_dataIn_W[35]
  PIN dyn0_dataIn_W[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 2496.000 1533.090 2500.000 ;
    END
  END dyn0_dataIn_W[36]
  PIN dyn0_dataIn_W[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2247.440 4.000 2248.040 ;
    END
  END dyn0_dataIn_W[37]
  PIN dyn0_dataIn_W[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END dyn0_dataIn_W[38]
  PIN dyn0_dataIn_W[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 4.000 ;
    END
  END dyn0_dataIn_W[39]
  PIN dyn0_dataIn_W[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 251.640 2500.000 252.240 ;
    END
  END dyn0_dataIn_W[3]
  PIN dyn0_dataIn_W[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END dyn0_dataIn_W[40]
  PIN dyn0_dataIn_W[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2179.440 4.000 2180.040 ;
    END
  END dyn0_dataIn_W[41]
  PIN dyn0_dataIn_W[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 299.240 2500.000 299.840 ;
    END
  END dyn0_dataIn_W[42]
  PIN dyn0_dataIn_W[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 4.000 1292.640 ;
    END
  END dyn0_dataIn_W[43]
  PIN dyn0_dataIn_W[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2125.040 4.000 2125.640 ;
    END
  END dyn0_dataIn_W[44]
  PIN dyn0_dataIn_W[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END dyn0_dataIn_W[45]
  PIN dyn0_dataIn_W[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 4.000 ;
    END
  END dyn0_dataIn_W[46]
  PIN dyn0_dataIn_W[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1139.040 2500.000 1139.640 ;
    END
  END dyn0_dataIn_W[47]
  PIN dyn0_dataIn_W[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END dyn0_dataIn_W[48]
  PIN dyn0_dataIn_W[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 0.000 1719.850 4.000 ;
    END
  END dyn0_dataIn_W[49]
  PIN dyn0_dataIn_W[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 2496.000 1867.970 2500.000 ;
    END
  END dyn0_dataIn_W[4]
  PIN dyn0_dataIn_W[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1445.040 2500.000 1445.640 ;
    END
  END dyn0_dataIn_W[50]
  PIN dyn0_dataIn_W[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 350.240 2500.000 350.840 ;
    END
  END dyn0_dataIn_W[51]
  PIN dyn0_dataIn_W[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1383.840 2500.000 1384.440 ;
    END
  END dyn0_dataIn_W[52]
  PIN dyn0_dataIn_W[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END dyn0_dataIn_W[53]
  PIN dyn0_dataIn_W[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.470 0.000 2347.750 4.000 ;
    END
  END dyn0_dataIn_W[54]
  PIN dyn0_dataIn_W[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2383.440 2500.000 2384.040 ;
    END
  END dyn0_dataIn_W[55]
  PIN dyn0_dataIn_W[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.870 0.000 2412.150 4.000 ;
    END
  END dyn0_dataIn_W[56]
  PIN dyn0_dataIn_W[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 2496.000 1787.470 2500.000 ;
    END
  END dyn0_dataIn_W[57]
  PIN dyn0_dataIn_W[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 2496.000 174.250 2500.000 ;
    END
  END dyn0_dataIn_W[58]
  PIN dyn0_dataIn_W[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END dyn0_dataIn_W[59]
  PIN dyn0_dataIn_W[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 717.440 2500.000 718.040 ;
    END
  END dyn0_dataIn_W[5]
  PIN dyn0_dataIn_W[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 0.000 1771.370 4.000 ;
    END
  END dyn0_dataIn_W[60]
  PIN dyn0_dataIn_W[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 601.840 2500.000 602.440 ;
    END
  END dyn0_dataIn_W[61]
  PIN dyn0_dataIn_W[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2152.240 4.000 2152.840 ;
    END
  END dyn0_dataIn_W[62]
  PIN dyn0_dataIn_W[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.240 4.000 1574.840 ;
    END
  END dyn0_dataIn_W[63]
  PIN dyn0_dataIn_W[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END dyn0_dataIn_W[6]
  PIN dyn0_dataIn_W[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 2496.000 715.210 2500.000 ;
    END
  END dyn0_dataIn_W[7]
  PIN dyn0_dataIn_W[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END dyn0_dataIn_W[8]
  PIN dyn0_dataIn_W[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1706.840 2500.000 1707.440 ;
    END
  END dyn0_dataIn_W[9]
  PIN dyn0_validIn_E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.570 2496.000 2363.850 2500.000 ;
    END
  END dyn0_validIn_E
  PIN dyn0_validIn_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2403.840 2500.000 2404.440 ;
    END
  END dyn0_validIn_N
  PIN dyn0_validIn_S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END dyn0_validIn_S
  PIN dyn0_validIn_W
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END dyn0_validIn_W
  PIN dyn0_yummyOut_E
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 0.000 1871.190 4.000 ;
    END
  END dyn0_yummyOut_E
  PIN dyn0_yummyOut_N
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END dyn0_yummyOut_N
  PIN dyn0_yummyOut_S
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 2496.000 1729.510 2500.000 ;
    END
  END dyn0_yummyOut_S
  PIN dyn0_yummyOut_W
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2006.040 2500.000 2006.640 ;
    END
  END dyn0_yummyOut_W
  PIN dyn1_dEo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 401.240 2500.000 401.840 ;
    END
  END dyn1_dEo[0]
  PIN dyn1_dEo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END dyn1_dEo[10]
  PIN dyn1_dEo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2478.640 4.000 2479.240 ;
    END
  END dyn1_dEo[11]
  PIN dyn1_dEo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END dyn1_dEo[12]
  PIN dyn1_dEo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2074.040 4.000 2074.640 ;
    END
  END dyn1_dEo[13]
  PIN dyn1_dEo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END dyn1_dEo[14]
  PIN dyn1_dEo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1853.040 4.000 1853.640 ;
    END
  END dyn1_dEo[15]
  PIN dyn1_dEo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END dyn1_dEo[16]
  PIN dyn1_dEo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1441.640 4.000 1442.240 ;
    END
  END dyn1_dEo[17]
  PIN dyn1_dEo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1105.040 2500.000 1105.640 ;
    END
  END dyn1_dEo[18]
  PIN dyn1_dEo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1264.840 2500.000 1265.440 ;
    END
  END dyn1_dEo[19]
  PIN dyn1_dEo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2172.640 4.000 2173.240 ;
    END
  END dyn1_dEo[1]
  PIN dyn1_dEo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END dyn1_dEo[20]
  PIN dyn1_dEo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 0.000 2241.490 4.000 ;
    END
  END dyn1_dEo[21]
  PIN dyn1_dEo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END dyn1_dEo[22]
  PIN dyn1_dEo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.430 2496.000 2405.710 2500.000 ;
    END
  END dyn1_dEo[23]
  PIN dyn1_dEo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1822.440 4.000 1823.040 ;
    END
  END dyn1_dEo[24]
  PIN dyn1_dEo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1373.640 4.000 1374.240 ;
    END
  END dyn1_dEo[25]
  PIN dyn1_dEo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END dyn1_dEo[26]
  PIN dyn1_dEo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END dyn1_dEo[27]
  PIN dyn1_dEo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.410 2496.000 2273.690 2500.000 ;
    END
  END dyn1_dEo[28]
  PIN dyn1_dEo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END dyn1_dEo[29]
  PIN dyn1_dEo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 2496.000 724.870 2500.000 ;
    END
  END dyn1_dEo[2]
  PIN dyn1_dEo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END dyn1_dEo[30]
  PIN dyn1_dEo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.770 0.000 2235.050 4.000 ;
    END
  END dyn1_dEo[31]
  PIN dyn1_dEo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END dyn1_dEo[32]
  PIN dyn1_dEo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 2496.000 1220.750 2500.000 ;
    END
  END dyn1_dEo[33]
  PIN dyn1_dEo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END dyn1_dEo[34]
  PIN dyn1_dEo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END dyn1_dEo[35]
  PIN dyn1_dEo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 2496.000 322.370 2500.000 ;
    END
  END dyn1_dEo[36]
  PIN dyn1_dEo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END dyn1_dEo[37]
  PIN dyn1_dEo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 2496.000 821.470 2500.000 ;
    END
  END dyn1_dEo[38]
  PIN dyn1_dEo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2043.440 4.000 2044.040 ;
    END
  END dyn1_dEo[39]
  PIN dyn1_dEo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END dyn1_dEo[3]
  PIN dyn1_dEo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 2496.000 956.710 2500.000 ;
    END
  END dyn1_dEo[40]
  PIN dyn1_dEo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 2496.000 895.530 2500.000 ;
    END
  END dyn1_dEo[41]
  PIN dyn1_dEo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1339.640 2500.000 1340.240 ;
    END
  END dyn1_dEo[42]
  PIN dyn1_dEo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END dyn1_dEo[43]
  PIN dyn1_dEo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 2496.000 1516.990 2500.000 ;
    END
  END dyn1_dEo[44]
  PIN dyn1_dEo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1482.440 2500.000 1483.040 ;
    END
  END dyn1_dEo[45]
  PIN dyn1_dEo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 547.440 2500.000 548.040 ;
    END
  END dyn1_dEo[46]
  PIN dyn1_dEo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END dyn1_dEo[47]
  PIN dyn1_dEo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END dyn1_dEo[48]
  PIN dyn1_dEo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2097.840 2500.000 2098.440 ;
    END
  END dyn1_dEo[49]
  PIN dyn1_dEo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END dyn1_dEo[4]
  PIN dyn1_dEo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END dyn1_dEo[50]
  PIN dyn1_dEo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1819.040 4.000 1819.640 ;
    END
  END dyn1_dEo[51]
  PIN dyn1_dEo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END dyn1_dEo[52]
  PIN dyn1_dEo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 0.000 1285.150 4.000 ;
    END
  END dyn1_dEo[53]
  PIN dyn1_dEo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.840 4.000 1520.440 ;
    END
  END dyn1_dEo[54]
  PIN dyn1_dEo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 2496.000 2086.930 2500.000 ;
    END
  END dyn1_dEo[55]
  PIN dyn1_dEo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1465.440 2500.000 1466.040 ;
    END
  END dyn1_dEo[56]
  PIN dyn1_dEo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 2496.000 1842.210 2500.000 ;
    END
  END dyn1_dEo[57]
  PIN dyn1_dEo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2196.440 4.000 2197.040 ;
    END
  END dyn1_dEo[58]
  PIN dyn1_dEo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 0.000 1581.390 4.000 ;
    END
  END dyn1_dEo[59]
  PIN dyn1_dEo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2121.640 4.000 2122.240 ;
    END
  END dyn1_dEo[5]
  PIN dyn1_dEo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END dyn1_dEo[60]
  PIN dyn1_dEo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 2496.000 937.390 2500.000 ;
    END
  END dyn1_dEo[61]
  PIN dyn1_dEo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END dyn1_dEo[62]
  PIN dyn1_dEo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 0.000 1922.710 4.000 ;
    END
  END dyn1_dEo[63]
  PIN dyn1_dEo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1815.640 4.000 1816.240 ;
    END
  END dyn1_dEo[6]
  PIN dyn1_dEo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 2496.000 106.630 2500.000 ;
    END
  END dyn1_dEo[7]
  PIN dyn1_dEo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END dyn1_dEo[8]
  PIN dyn1_dEo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.790 2496.000 1723.070 2500.000 ;
    END
  END dyn1_dEo[9]
  PIN dyn1_dEo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END dyn1_dEo_valid
  PIN dyn1_dEo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END dyn1_dEo_yummy
  PIN dyn1_dNo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END dyn1_dNo[0]
  PIN dyn1_dNo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END dyn1_dNo[10]
  PIN dyn1_dNo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 2496.000 1259.390 2500.000 ;
    END
  END dyn1_dNo[11]
  PIN dyn1_dNo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END dyn1_dNo[12]
  PIN dyn1_dNo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END dyn1_dNo[13]
  PIN dyn1_dNo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 214.240 2500.000 214.840 ;
    END
  END dyn1_dNo[14]
  PIN dyn1_dNo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1186.640 4.000 1187.240 ;
    END
  END dyn1_dNo[15]
  PIN dyn1_dNo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2145.440 2500.000 2146.040 ;
    END
  END dyn1_dNo[16]
  PIN dyn1_dNo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END dyn1_dNo[17]
  PIN dyn1_dNo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2407.240 2500.000 2407.840 ;
    END
  END dyn1_dNo[18]
  PIN dyn1_dNo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END dyn1_dNo[19]
  PIN dyn1_dNo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2213.440 4.000 2214.040 ;
    END
  END dyn1_dNo[1]
  PIN dyn1_dNo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 2496.000 905.190 2500.000 ;
    END
  END dyn1_dNo[20]
  PIN dyn1_dNo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 2496.000 856.890 2500.000 ;
    END
  END dyn1_dNo[21]
  PIN dyn1_dNo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 2496.000 1088.730 2500.000 ;
    END
  END dyn1_dNo[22]
  PIN dyn1_dNo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END dyn1_dNo[23]
  PIN dyn1_dNo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 870.440 2500.000 871.040 ;
    END
  END dyn1_dNo[24]
  PIN dyn1_dNo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1581.040 4.000 1581.640 ;
    END
  END dyn1_dNo[25]
  PIN dyn1_dNo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END dyn1_dNo[26]
  PIN dyn1_dNo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END dyn1_dNo[27]
  PIN dyn1_dNo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 2496.000 2125.570 2500.000 ;
    END
  END dyn1_dNo[28]
  PIN dyn1_dNo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END dyn1_dNo[29]
  PIN dyn1_dNo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2478.640 2500.000 2479.240 ;
    END
  END dyn1_dNo[2]
  PIN dyn1_dNo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2339.240 4.000 2339.840 ;
    END
  END dyn1_dNo[30]
  PIN dyn1_dNo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1302.240 2500.000 1302.840 ;
    END
  END dyn1_dNo[31]
  PIN dyn1_dNo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 0.000 1748.830 4.000 ;
    END
  END dyn1_dNo[32]
  PIN dyn1_dNo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2298.440 4.000 2299.040 ;
    END
  END dyn1_dNo[33]
  PIN dyn1_dNo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 826.240 2500.000 826.840 ;
    END
  END dyn1_dNo[34]
  PIN dyn1_dNo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1642.240 2500.000 1642.840 ;
    END
  END dyn1_dNo[35]
  PIN dyn1_dNo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 2496.000 138.830 2500.000 ;
    END
  END dyn1_dNo[36]
  PIN dyn1_dNo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.490 0.000 2157.770 4.000 ;
    END
  END dyn1_dNo[37]
  PIN dyn1_dNo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1672.840 2500.000 1673.440 ;
    END
  END dyn1_dNo[38]
  PIN dyn1_dNo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2053.640 4.000 2054.240 ;
    END
  END dyn1_dNo[39]
  PIN dyn1_dNo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1207.040 2500.000 1207.640 ;
    END
  END dyn1_dNo[3]
  PIN dyn1_dNo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1448.440 2500.000 1449.040 ;
    END
  END dyn1_dNo[40]
  PIN dyn1_dNo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.150 2496.000 2006.430 2500.000 ;
    END
  END dyn1_dNo[41]
  PIN dyn1_dNo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690 0.000 2350.970 4.000 ;
    END
  END dyn1_dNo[42]
  PIN dyn1_dNo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 2496.000 950.270 2500.000 ;
    END
  END dyn1_dNo[43]
  PIN dyn1_dNo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2308.830 2496.000 2309.110 2500.000 ;
    END
  END dyn1_dNo[44]
  PIN dyn1_dNo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2475.240 4.000 2475.840 ;
    END
  END dyn1_dNo[45]
  PIN dyn1_dNo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 2496.000 1137.030 2500.000 ;
    END
  END dyn1_dNo[46]
  PIN dyn1_dNo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1880.240 2500.000 1880.840 ;
    END
  END dyn1_dNo[47]
  PIN dyn1_dNo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2240.640 2500.000 2241.240 ;
    END
  END dyn1_dNo[48]
  PIN dyn1_dNo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END dyn1_dNo[49]
  PIN dyn1_dNo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END dyn1_dNo[4]
  PIN dyn1_dNo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 224.440 2500.000 225.040 ;
    END
  END dyn1_dNo[50]
  PIN dyn1_dNo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END dyn1_dNo[51]
  PIN dyn1_dNo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 574.640 2500.000 575.240 ;
    END
  END dyn1_dNo[52]
  PIN dyn1_dNo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END dyn1_dNo[53]
  PIN dyn1_dNo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1883.640 4.000 1884.240 ;
    END
  END dyn1_dNo[54]
  PIN dyn1_dNo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END dyn1_dNo[55]
  PIN dyn1_dNo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 489.640 2500.000 490.240 ;
    END
  END dyn1_dNo[56]
  PIN dyn1_dNo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 2496.000 621.830 2500.000 ;
    END
  END dyn1_dNo[57]
  PIN dyn1_dNo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1774.840 4.000 1775.440 ;
    END
  END dyn1_dNo[58]
  PIN dyn1_dNo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 2496.000 631.490 2500.000 ;
    END
  END dyn1_dNo[59]
  PIN dyn1_dNo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.840 4.000 1554.440 ;
    END
  END dyn1_dNo[5]
  PIN dyn1_dNo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 894.240 2500.000 894.840 ;
    END
  END dyn1_dNo[60]
  PIN dyn1_dNo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2393.640 4.000 2394.240 ;
    END
  END dyn1_dNo[61]
  PIN dyn1_dNo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END dyn1_dNo[62]
  PIN dyn1_dNo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2210.040 4.000 2210.640 ;
    END
  END dyn1_dNo[63]
  PIN dyn1_dNo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1400.840 2500.000 1401.440 ;
    END
  END dyn1_dNo[6]
  PIN dyn1_dNo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END dyn1_dNo[7]
  PIN dyn1_dNo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 2496.000 1488.010 2500.000 ;
    END
  END dyn1_dNo[8]
  PIN dyn1_dNo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END dyn1_dNo[9]
  PIN dyn1_dNo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 2496.000 1719.850 2500.000 ;
    END
  END dyn1_dNo_valid
  PIN dyn1_dNo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 4.000 ;
    END
  END dyn1_dNo_yummy
  PIN dyn1_dSo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 2496.000 1021.110 2500.000 ;
    END
  END dyn1_dSo[0]
  PIN dyn1_dSo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.150 0.000 2167.430 4.000 ;
    END
  END dyn1_dSo[10]
  PIN dyn1_dSo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END dyn1_dSo[11]
  PIN dyn1_dSo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 2496.000 116.290 2500.000 ;
    END
  END dyn1_dSo[12]
  PIN dyn1_dSo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END dyn1_dSo[13]
  PIN dyn1_dSo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END dyn1_dSo[14]
  PIN dyn1_dSo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 2496.000 592.850 2500.000 ;
    END
  END dyn1_dSo[15]
  PIN dyn1_dSo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END dyn1_dSo[16]
  PIN dyn1_dSo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 404.640 2500.000 405.240 ;
    END
  END dyn1_dSo[17]
  PIN dyn1_dSo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 2496.000 744.190 2500.000 ;
    END
  END dyn1_dSo[18]
  PIN dyn1_dSo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END dyn1_dSo[19]
  PIN dyn1_dSo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 2496.000 692.670 2500.000 ;
    END
  END dyn1_dSo[1]
  PIN dyn1_dSo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END dyn1_dSo[20]
  PIN dyn1_dSo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1587.840 4.000 1588.440 ;
    END
  END dyn1_dSo[21]
  PIN dyn1_dSo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1132.240 2500.000 1132.840 ;
    END
  END dyn1_dSo[22]
  PIN dyn1_dSo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.030 2496.000 2180.310 2500.000 ;
    END
  END dyn1_dSo[23]
  PIN dyn1_dSo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END dyn1_dSo[24]
  PIN dyn1_dSo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1941.440 2500.000 1942.040 ;
    END
  END dyn1_dSo[25]
  PIN dyn1_dSo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 0.000 2270.470 4.000 ;
    END
  END dyn1_dSo[26]
  PIN dyn1_dSo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2244.040 4.000 2244.640 ;
    END
  END dyn1_dSo[27]
  PIN dyn1_dSo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 2496.000 1410.730 2500.000 ;
    END
  END dyn1_dSo[28]
  PIN dyn1_dSo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 2496.000 914.850 2500.000 ;
    END
  END dyn1_dSo[29]
  PIN dyn1_dSo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1890.440 2500.000 1891.040 ;
    END
  END dyn1_dSo[2]
  PIN dyn1_dSo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1298.840 2500.000 1299.440 ;
    END
  END dyn1_dSo[30]
  PIN dyn1_dSo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 537.240 2500.000 537.840 ;
    END
  END dyn1_dSo[31]
  PIN dyn1_dSo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END dyn1_dSo[32]
  PIN dyn1_dSo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 2496.000 824.690 2500.000 ;
    END
  END dyn1_dSo[33]
  PIN dyn1_dSo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2431.040 4.000 2431.640 ;
    END
  END dyn1_dSo[34]
  PIN dyn1_dSo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1411.040 2500.000 1411.640 ;
    END
  END dyn1_dSo[35]
  PIN dyn1_dSo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END dyn1_dSo[36]
  PIN dyn1_dSo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END dyn1_dSo[37]
  PIN dyn1_dSo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 741.240 2500.000 741.840 ;
    END
  END dyn1_dSo[38]
  PIN dyn1_dSo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END dyn1_dSo[39]
  PIN dyn1_dSo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 2496.000 29.350 2500.000 ;
    END
  END dyn1_dSo[3]
  PIN dyn1_dSo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1944.840 2500.000 1945.440 ;
    END
  END dyn1_dSo[40]
  PIN dyn1_dSo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1438.240 2500.000 1438.840 ;
    END
  END dyn1_dSo[41]
  PIN dyn1_dSo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END dyn1_dSo[42]
  PIN dyn1_dSo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.490 2496.000 1996.770 2500.000 ;
    END
  END dyn1_dSo[43]
  PIN dyn1_dSo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 2496.000 473.710 2500.000 ;
    END
  END dyn1_dSo[44]
  PIN dyn1_dSo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1506.240 4.000 1506.840 ;
    END
  END dyn1_dSo[45]
  PIN dyn1_dSo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1023.440 2500.000 1024.040 ;
    END
  END dyn1_dSo[46]
  PIN dyn1_dSo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 523.640 2500.000 524.240 ;
    END
  END dyn1_dSo[47]
  PIN dyn1_dSo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 435.240 2500.000 435.840 ;
    END
  END dyn1_dSo[48]
  PIN dyn1_dSo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2295.040 4.000 2295.640 ;
    END
  END dyn1_dSo[49]
  PIN dyn1_dSo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.240 4.000 1336.840 ;
    END
  END dyn1_dSo[4]
  PIN dyn1_dSo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 122.440 2500.000 123.040 ;
    END
  END dyn1_dSo[50]
  PIN dyn1_dSo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1149.240 2500.000 1149.840 ;
    END
  END dyn1_dSo[51]
  PIN dyn1_dSo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END dyn1_dSo[52]
  PIN dyn1_dSo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.510 2496.000 2289.790 2500.000 ;
    END
  END dyn1_dSo[53]
  PIN dyn1_dSo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END dyn1_dSo[54]
  PIN dyn1_dSo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END dyn1_dSo[55]
  PIN dyn1_dSo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2410.640 2500.000 2411.240 ;
    END
  END dyn1_dSo[56]
  PIN dyn1_dSo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2444.640 4.000 2445.240 ;
    END
  END dyn1_dSo[57]
  PIN dyn1_dSo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2023.040 2500.000 2023.640 ;
    END
  END dyn1_dSo[58]
  PIN dyn1_dSo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2284.840 4.000 2285.440 ;
    END
  END dyn1_dSo[59]
  PIN dyn1_dSo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END dyn1_dSo[5]
  PIN dyn1_dSo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END dyn1_dSo[60]
  PIN dyn1_dSo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2376.640 4.000 2377.240 ;
    END
  END dyn1_dSo[61]
  PIN dyn1_dSo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1570.840 2500.000 1571.440 ;
    END
  END dyn1_dSo[62]
  PIN dyn1_dSo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END dyn1_dSo[63]
  PIN dyn1_dSo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 2496.000 747.410 2500.000 ;
    END
  END dyn1_dSo[6]
  PIN dyn1_dSo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 2496.000 766.730 2500.000 ;
    END
  END dyn1_dSo[7]
  PIN dyn1_dSo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END dyn1_dSo[8]
  PIN dyn1_dSo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1978.840 2500.000 1979.440 ;
    END
  END dyn1_dSo[9]
  PIN dyn1_dSo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1856.440 2500.000 1857.040 ;
    END
  END dyn1_dSo_valid
  PIN dyn1_dSo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END dyn1_dSo_yummy
  PIN dyn1_dWo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END dyn1_dWo[0]
  PIN dyn1_dWo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END dyn1_dWo[10]
  PIN dyn1_dWo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.570 0.000 2041.850 4.000 ;
    END
  END dyn1_dWo[11]
  PIN dyn1_dWo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END dyn1_dWo[12]
  PIN dyn1_dWo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END dyn1_dWo[13]
  PIN dyn1_dWo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.070 0.000 2444.350 4.000 ;
    END
  END dyn1_dWo[14]
  PIN dyn1_dWo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 758.240 2500.000 758.840 ;
    END
  END dyn1_dWo[15]
  PIN dyn1_dWo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1863.240 4.000 1863.840 ;
    END
  END dyn1_dWo[16]
  PIN dyn1_dWo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1210.440 4.000 1211.040 ;
    END
  END dyn1_dWo[17]
  PIN dyn1_dWo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END dyn1_dWo[18]
  PIN dyn1_dWo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1574.240 2500.000 1574.840 ;
    END
  END dyn1_dWo[19]
  PIN dyn1_dWo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.530 2496.000 2260.810 2500.000 ;
    END
  END dyn1_dWo[1]
  PIN dyn1_dWo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 2496.000 293.390 2500.000 ;
    END
  END dyn1_dWo[20]
  PIN dyn1_dWo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.850 2496.000 2280.130 2500.000 ;
    END
  END dyn1_dWo[21]
  PIN dyn1_dWo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.730 0.000 1971.010 4.000 ;
    END
  END dyn1_dWo[22]
  PIN dyn1_dWo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 2496.000 795.710 2500.000 ;
    END
  END dyn1_dWo[23]
  PIN dyn1_dWo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 911.240 2500.000 911.840 ;
    END
  END dyn1_dWo[24]
  PIN dyn1_dWo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 2496.000 1101.610 2500.000 ;
    END
  END dyn1_dWo[25]
  PIN dyn1_dWo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END dyn1_dWo[26]
  PIN dyn1_dWo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END dyn1_dWo[27]
  PIN dyn1_dWo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 2496.000 1603.930 2500.000 ;
    END
  END dyn1_dWo[28]
  PIN dyn1_dWo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.190 2496.000 1626.470 2500.000 ;
    END
  END dyn1_dWo[29]
  PIN dyn1_dWo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END dyn1_dWo[2]
  PIN dyn1_dWo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 792.240 2500.000 792.840 ;
    END
  END dyn1_dWo[30]
  PIN dyn1_dWo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END dyn1_dWo[31]
  PIN dyn1_dWo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END dyn1_dWo[32]
  PIN dyn1_dWo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 2496.000 1236.850 2500.000 ;
    END
  END dyn1_dWo[33]
  PIN dyn1_dWo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END dyn1_dWo[34]
  PIN dyn1_dWo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2267.840 2500.000 2268.440 ;
    END
  END dyn1_dWo[35]
  PIN dyn1_dWo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.670 2496.000 2379.950 2500.000 ;
    END
  END dyn1_dWo[36]
  PIN dyn1_dWo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 2496.000 1942.030 2500.000 ;
    END
  END dyn1_dWo[37]
  PIN dyn1_dWo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2070.640 2500.000 2071.240 ;
    END
  END dyn1_dWo[38]
  PIN dyn1_dWo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 2496.000 1413.950 2500.000 ;
    END
  END dyn1_dWo[39]
  PIN dyn1_dWo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END dyn1_dWo[3]
  PIN dyn1_dWo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 2496.000 470.490 2500.000 ;
    END
  END dyn1_dWo[40]
  PIN dyn1_dWo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.930 0.000 2003.210 4.000 ;
    END
  END dyn1_dWo[41]
  PIN dyn1_dWo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.250 2496.000 2022.530 2500.000 ;
    END
  END dyn1_dWo[42]
  PIN dyn1_dWo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END dyn1_dWo[43]
  PIN dyn1_dWo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 244.840 2500.000 245.440 ;
    END
  END dyn1_dWo[44]
  PIN dyn1_dWo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 2496.000 1188.550 2500.000 ;
    END
  END dyn1_dWo[45]
  PIN dyn1_dWo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END dyn1_dWo[46]
  PIN dyn1_dWo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END dyn1_dWo[47]
  PIN dyn1_dWo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END dyn1_dWo[48]
  PIN dyn1_dWo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.370 0.000 2170.650 4.000 ;
    END
  END dyn1_dWo[49]
  PIN dyn1_dWo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 754.840 2500.000 755.440 ;
    END
  END dyn1_dWo[4]
  PIN dyn1_dWo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.730 2496.000 2454.010 2500.000 ;
    END
  END dyn1_dWo[50]
  PIN dyn1_dWo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 2496.000 216.110 2500.000 ;
    END
  END dyn1_dWo[51]
  PIN dyn1_dWo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END dyn1_dWo[52]
  PIN dyn1_dWo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 2496.000 200.010 2500.000 ;
    END
  END dyn1_dWo[53]
  PIN dyn1_dWo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2006.040 4.000 2006.640 ;
    END
  END dyn1_dWo[54]
  PIN dyn1_dWo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2223.640 4.000 2224.240 ;
    END
  END dyn1_dWo[55]
  PIN dyn1_dWo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 2496.000 1452.590 2500.000 ;
    END
  END dyn1_dWo[56]
  PIN dyn1_dWo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1846.240 4.000 1846.840 ;
    END
  END dyn1_dWo[57]
  PIN dyn1_dWo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 2496.000 1752.050 2500.000 ;
    END
  END dyn1_dWo[58]
  PIN dyn1_dWo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2023.040 4.000 2023.640 ;
    END
  END dyn1_dWo[59]
  PIN dyn1_dWo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END dyn1_dWo[5]
  PIN dyn1_dWo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2155.640 4.000 2156.240 ;
    END
  END dyn1_dWo[60]
  PIN dyn1_dWo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 2496.000 943.830 2500.000 ;
    END
  END dyn1_dWo[61]
  PIN dyn1_dWo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 4.000 ;
    END
  END dyn1_dWo[62]
  PIN dyn1_dWo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.090 2496.000 2254.370 2500.000 ;
    END
  END dyn1_dWo[63]
  PIN dyn1_dWo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END dyn1_dWo[6]
  PIN dyn1_dWo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 2496.000 1201.430 2500.000 ;
    END
  END dyn1_dWo[7]
  PIN dyn1_dWo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 0.000 1169.230 4.000 ;
    END
  END dyn1_dWo[8]
  PIN dyn1_dWo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1897.240 4.000 1897.840 ;
    END
  END dyn1_dWo[9]
  PIN dyn1_dWo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END dyn1_dWo_valid
  PIN dyn1_dWo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1485.840 2500.000 1486.440 ;
    END
  END dyn1_dWo_yummy
  PIN dyn1_dataIn_E[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1125.440 4.000 1126.040 ;
    END
  END dyn1_dataIn_E[0]
  PIN dyn1_dataIn_E[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 2496.000 1864.750 2500.000 ;
    END
  END dyn1_dataIn_E[10]
  PIN dyn1_dataIn_E[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 928.240 2500.000 928.840 ;
    END
  END dyn1_dataIn_E[11]
  PIN dyn1_dataIn_E[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 0.000 1629.690 4.000 ;
    END
  END dyn1_dataIn_E[12]
  PIN dyn1_dataIn_E[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.910 0.000 2193.190 4.000 ;
    END
  END dyn1_dataIn_E[13]
  PIN dyn1_dataIn_E[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END dyn1_dataIn_E[14]
  PIN dyn1_dataIn_E[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 0.000 1810.010 4.000 ;
    END
  END dyn1_dataIn_E[15]
  PIN dyn1_dataIn_E[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1366.840 2500.000 1367.440 ;
    END
  END dyn1_dataIn_E[16]
  PIN dyn1_dataIn_E[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1428.040 2500.000 1428.640 ;
    END
  END dyn1_dataIn_E[17]
  PIN dyn1_dataIn_E[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END dyn1_dataIn_E[18]
  PIN dyn1_dataIn_E[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.130 0.000 2035.410 4.000 ;
    END
  END dyn1_dataIn_E[19]
  PIN dyn1_dataIn_E[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 132.640 2500.000 133.240 ;
    END
  END dyn1_dataIn_E[1]
  PIN dyn1_dataIn_E[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 2496.000 241.870 2500.000 ;
    END
  END dyn1_dataIn_E[20]
  PIN dyn1_dataIn_E[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1992.440 2500.000 1993.040 ;
    END
  END dyn1_dataIn_E[21]
  PIN dyn1_dataIn_E[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END dyn1_dataIn_E[22]
  PIN dyn1_dataIn_E[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 2496.000 683.010 2500.000 ;
    END
  END dyn1_dataIn_E[23]
  PIN dyn1_dataIn_E[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.330 0.000 1101.610 4.000 ;
    END
  END dyn1_dataIn_E[24]
  PIN dyn1_dataIn_E[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 0.000 2312.330 4.000 ;
    END
  END dyn1_dataIn_E[25]
  PIN dyn1_dataIn_E[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 642.640 2500.000 643.240 ;
    END
  END dyn1_dataIn_E[26]
  PIN dyn1_dataIn_E[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END dyn1_dataIn_E[27]
  PIN dyn1_dataIn_E[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1921.040 2500.000 1921.640 ;
    END
  END dyn1_dataIn_E[28]
  PIN dyn1_dataIn_E[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END dyn1_dataIn_E[29]
  PIN dyn1_dataIn_E[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END dyn1_dataIn_E[2]
  PIN dyn1_dataIn_E[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 2496.000 763.510 2500.000 ;
    END
  END dyn1_dataIn_E[30]
  PIN dyn1_dataIn_E[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2373.240 2500.000 2373.840 ;
    END
  END dyn1_dataIn_E[31]
  PIN dyn1_dataIn_E[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1924.440 2500.000 1925.040 ;
    END
  END dyn1_dataIn_E[32]
  PIN dyn1_dataIn_E[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.490 0.000 2318.770 4.000 ;
    END
  END dyn1_dataIn_E[33]
  PIN dyn1_dataIn_E[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2329.040 4.000 2329.640 ;
    END
  END dyn1_dataIn_E[34]
  PIN dyn1_dataIn_E[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 4.000 ;
    END
  END dyn1_dataIn_E[35]
  PIN dyn1_dataIn_E[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 2496.000 898.750 2500.000 ;
    END
  END dyn1_dataIn_E[36]
  PIN dyn1_dataIn_E[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1237.640 2500.000 1238.240 ;
    END
  END dyn1_dataIn_E[37]
  PIN dyn1_dataIn_E[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END dyn1_dataIn_E[38]
  PIN dyn1_dataIn_E[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 2496.000 1388.190 2500.000 ;
    END
  END dyn1_dataIn_E[39]
  PIN dyn1_dataIn_E[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END dyn1_dataIn_E[3]
  PIN dyn1_dataIn_E[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.010 0.000 2370.290 4.000 ;
    END
  END dyn1_dataIn_E[40]
  PIN dyn1_dataIn_E[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END dyn1_dataIn_E[41]
  PIN dyn1_dataIn_E[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 2496.000 547.770 2500.000 ;
    END
  END dyn1_dataIn_E[42]
  PIN dyn1_dataIn_E[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 513.440 2500.000 514.040 ;
    END
  END dyn1_dataIn_E[43]
  PIN dyn1_dataIn_E[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 2496.000 1764.930 2500.000 ;
    END
  END dyn1_dataIn_E[44]
  PIN dyn1_dataIn_E[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1649.040 2500.000 1649.640 ;
    END
  END dyn1_dataIn_E[45]
  PIN dyn1_dataIn_E[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 2496.000 599.290 2500.000 ;
    END
  END dyn1_dataIn_E[46]
  PIN dyn1_dataIn_E[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END dyn1_dataIn_E[47]
  PIN dyn1_dataIn_E[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1322.640 2500.000 1323.240 ;
    END
  END dyn1_dataIn_E[48]
  PIN dyn1_dataIn_E[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1312.440 2500.000 1313.040 ;
    END
  END dyn1_dataIn_E[49]
  PIN dyn1_dataIn_E[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 4.000 2455.440 ;
    END
  END dyn1_dataIn_E[4]
  PIN dyn1_dataIn_E[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.690 0.000 2189.970 4.000 ;
    END
  END dyn1_dataIn_E[50]
  PIN dyn1_dataIn_E[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 0.000 1687.650 4.000 ;
    END
  END dyn1_dataIn_E[51]
  PIN dyn1_dataIn_E[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END dyn1_dataIn_E[52]
  PIN dyn1_dataIn_E[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END dyn1_dataIn_E[53]
  PIN dyn1_dataIn_E[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 0.000 1362.430 4.000 ;
    END
  END dyn1_dataIn_E[54]
  PIN dyn1_dataIn_E[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.050 0.000 2473.330 4.000 ;
    END
  END dyn1_dataIn_E[55]
  PIN dyn1_dataIn_E[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END dyn1_dataIn_E[56]
  PIN dyn1_dataIn_E[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END dyn1_dataIn_E[57]
  PIN dyn1_dataIn_E[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END dyn1_dataIn_E[58]
  PIN dyn1_dataIn_E[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END dyn1_dataIn_E[59]
  PIN dyn1_dataIn_E[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 2496.000 679.790 2500.000 ;
    END
  END dyn1_dataIn_E[5]
  PIN dyn1_dataIn_E[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 591.640 2500.000 592.240 ;
    END
  END dyn1_dataIn_E[60]
  PIN dyn1_dataIn_E[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 2496.000 982.470 2500.000 ;
    END
  END dyn1_dataIn_E[61]
  PIN dyn1_dataIn_E[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 2496.000 1761.710 2500.000 ;
    END
  END dyn1_dataIn_E[62]
  PIN dyn1_dataIn_E[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END dyn1_dataIn_E[63]
  PIN dyn1_dataIn_E[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.770 2496.000 2074.050 2500.000 ;
    END
  END dyn1_dataIn_E[6]
  PIN dyn1_dataIn_E[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END dyn1_dataIn_E[7]
  PIN dyn1_dataIn_E[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END dyn1_dataIn_E[8]
  PIN dyn1_dataIn_E[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 2496.000 1378.530 2500.000 ;
    END
  END dyn1_dataIn_E[9]
  PIN dyn1_dataIn_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END dyn1_dataIn_N[0]
  PIN dyn1_dataIn_N[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1166.240 2500.000 1166.840 ;
    END
  END dyn1_dataIn_N[10]
  PIN dyn1_dataIn_N[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2335.840 4.000 2336.440 ;
    END
  END dyn1_dataIn_N[11]
  PIN dyn1_dataIn_N[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END dyn1_dataIn_N[12]
  PIN dyn1_dataIn_N[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1033.640 2500.000 1034.240 ;
    END
  END dyn1_dataIn_N[13]
  PIN dyn1_dataIn_N[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END dyn1_dataIn_N[14]
  PIN dyn1_dataIn_N[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2346.040 2500.000 2346.640 ;
    END
  END dyn1_dataIn_N[15]
  PIN dyn1_dataIn_N[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 2496.000 1230.410 2500.000 ;
    END
  END dyn1_dataIn_N[16]
  PIN dyn1_dataIn_N[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END dyn1_dataIn_N[17]
  PIN dyn1_dataIn_N[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END dyn1_dataIn_N[18]
  PIN dyn1_dataIn_N[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1934.640 2500.000 1935.240 ;
    END
  END dyn1_dataIn_N[19]
  PIN dyn1_dataIn_N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END dyn1_dataIn_N[1]
  PIN dyn1_dataIn_N[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 2496.000 1826.110 2500.000 ;
    END
  END dyn1_dataIn_N[20]
  PIN dyn1_dataIn_N[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2315.440 4.000 2316.040 ;
    END
  END dyn1_dataIn_N[21]
  PIN dyn1_dataIn_N[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1387.240 2500.000 1387.840 ;
    END
  END dyn1_dataIn_N[22]
  PIN dyn1_dataIn_N[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1458.640 2500.000 1459.240 ;
    END
  END dyn1_dataIn_N[23]
  PIN dyn1_dataIn_N[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1081.240 2500.000 1081.840 ;
    END
  END dyn1_dataIn_N[24]
  PIN dyn1_dataIn_N[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1502.840 2500.000 1503.440 ;
    END
  END dyn1_dataIn_N[25]
  PIN dyn1_dataIn_N[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 2496.000 270.850 2500.000 ;
    END
  END dyn1_dataIn_N[26]
  PIN dyn1_dataIn_N[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END dyn1_dataIn_N[27]
  PIN dyn1_dataIn_N[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END dyn1_dataIn_N[28]
  PIN dyn1_dataIn_N[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.970 0.000 1784.250 4.000 ;
    END
  END dyn1_dataIn_N[29]
  PIN dyn1_dataIn_N[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 2496.000 947.050 2500.000 ;
    END
  END dyn1_dataIn_N[2]
  PIN dyn1_dataIn_N[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END dyn1_dataIn_N[30]
  PIN dyn1_dataIn_N[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.630 2496.000 2437.910 2500.000 ;
    END
  END dyn1_dataIn_N[31]
  PIN dyn1_dataIn_N[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.410 0.000 2434.690 4.000 ;
    END
  END dyn1_dataIn_N[32]
  PIN dyn1_dataIn_N[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 802.440 2500.000 803.040 ;
    END
  END dyn1_dataIn_N[33]
  PIN dyn1_dataIn_N[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END dyn1_dataIn_N[34]
  PIN dyn1_dataIn_N[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.950 2496.000 1974.230 2500.000 ;
    END
  END dyn1_dataIn_N[35]
  PIN dyn1_dataIn_N[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 527.040 2500.000 527.640 ;
    END
  END dyn1_dataIn_N[36]
  PIN dyn1_dataIn_N[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END dyn1_dataIn_N[37]
  PIN dyn1_dataIn_N[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1499.440 2500.000 1500.040 ;
    END
  END dyn1_dataIn_N[38]
  PIN dyn1_dataIn_N[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 904.440 2500.000 905.040 ;
    END
  END dyn1_dataIn_N[39]
  PIN dyn1_dataIn_N[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 2496.000 274.070 2500.000 ;
    END
  END dyn1_dataIn_N[3]
  PIN dyn1_dataIn_N[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 2496.000 2119.130 2500.000 ;
    END
  END dyn1_dataIn_N[40]
  PIN dyn1_dataIn_N[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.430 0.000 2405.710 4.000 ;
    END
  END dyn1_dataIn_N[41]
  PIN dyn1_dataIn_N[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END dyn1_dataIn_N[42]
  PIN dyn1_dataIn_N[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END dyn1_dataIn_N[43]
  PIN dyn1_dataIn_N[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1836.040 4.000 1836.640 ;
    END
  END dyn1_dataIn_N[44]
  PIN dyn1_dataIn_N[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 2496.000 389.990 2500.000 ;
    END
  END dyn1_dataIn_N[45]
  PIN dyn1_dataIn_N[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 2496.000 1397.850 2500.000 ;
    END
  END dyn1_dataIn_N[46]
  PIN dyn1_dataIn_N[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END dyn1_dataIn_N[47]
  PIN dyn1_dataIn_N[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END dyn1_dataIn_N[48]
  PIN dyn1_dataIn_N[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END dyn1_dataIn_N[49]
  PIN dyn1_dataIn_N[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 2496.000 1658.670 2500.000 ;
    END
  END dyn1_dataIn_N[4]
  PIN dyn1_dataIn_N[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END dyn1_dataIn_N[50]
  PIN dyn1_dataIn_N[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2431.040 2500.000 2431.640 ;
    END
  END dyn1_dataIn_N[51]
  PIN dyn1_dataIn_N[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 23.840 2500.000 24.440 ;
    END
  END dyn1_dataIn_N[52]
  PIN dyn1_dataIn_N[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1506.240 2500.000 1506.840 ;
    END
  END dyn1_dataIn_N[53]
  PIN dyn1_dataIn_N[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2019.640 2500.000 2020.240 ;
    END
  END dyn1_dataIn_N[54]
  PIN dyn1_dataIn_N[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 156.440 2500.000 157.040 ;
    END
  END dyn1_dataIn_N[55]
  PIN dyn1_dataIn_N[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1676.240 2500.000 1676.840 ;
    END
  END dyn1_dataIn_N[56]
  PIN dyn1_dataIn_N[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 0.000 1243.290 4.000 ;
    END
  END dyn1_dataIn_N[57]
  PIN dyn1_dataIn_N[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 2496.000 283.730 2500.000 ;
    END
  END dyn1_dataIn_N[58]
  PIN dyn1_dataIn_N[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 2496.000 1813.230 2500.000 ;
    END
  END dyn1_dataIn_N[59]
  PIN dyn1_dataIn_N[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END dyn1_dataIn_N[5]
  PIN dyn1_dataIn_N[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1887.040 4.000 1887.640 ;
    END
  END dyn1_dataIn_N[60]
  PIN dyn1_dataIn_N[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 2496.000 1800.350 2500.000 ;
    END
  END dyn1_dataIn_N[61]
  PIN dyn1_dataIn_N[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 2496.000 402.870 2500.000 ;
    END
  END dyn1_dataIn_N[62]
  PIN dyn1_dataIn_N[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 2496.000 699.110 2500.000 ;
    END
  END dyn1_dataIn_N[63]
  PIN dyn1_dataIn_N[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.430 2496.000 2083.710 2500.000 ;
    END
  END dyn1_dataIn_N[6]
  PIN dyn1_dataIn_N[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.570 2496.000 2202.850 2500.000 ;
    END
  END dyn1_dataIn_N[7]
  PIN dyn1_dataIn_N[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1162.840 2500.000 1163.440 ;
    END
  END dyn1_dataIn_N[8]
  PIN dyn1_dataIn_N[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 0.000 1507.330 4.000 ;
    END
  END dyn1_dataIn_N[9]
  PIN dyn1_dataIn_S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 115.640 2500.000 116.240 ;
    END
  END dyn1_dataIn_S[0]
  PIN dyn1_dataIn_S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END dyn1_dataIn_S[10]
  PIN dyn1_dataIn_S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 663.040 2500.000 663.640 ;
    END
  END dyn1_dataIn_S[11]
  PIN dyn1_dataIn_S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 2496.000 248.310 2500.000 ;
    END
  END dyn1_dataIn_S[12]
  PIN dyn1_dataIn_S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.270 0.000 2476.550 4.000 ;
    END
  END dyn1_dataIn_S[13]
  PIN dyn1_dataIn_S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 567.840 2500.000 568.440 ;
    END
  END dyn1_dataIn_S[14]
  PIN dyn1_dataIn_S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2363.040 4.000 2363.640 ;
    END
  END dyn1_dataIn_S[15]
  PIN dyn1_dataIn_S[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 2496.000 737.750 2500.000 ;
    END
  END dyn1_dataIn_S[16]
  PIN dyn1_dataIn_S[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END dyn1_dataIn_S[17]
  PIN dyn1_dataIn_S[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1540.240 4.000 1540.840 ;
    END
  END dyn1_dataIn_S[18]
  PIN dyn1_dataIn_S[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 941.840 2500.000 942.440 ;
    END
  END dyn1_dataIn_S[19]
  PIN dyn1_dataIn_S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END dyn1_dataIn_S[1]
  PIN dyn1_dataIn_S[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 0.000 1800.350 4.000 ;
    END
  END dyn1_dataIn_S[20]
  PIN dyn1_dataIn_S[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 2496.000 1893.730 2500.000 ;
    END
  END dyn1_dataIn_S[21]
  PIN dyn1_dataIn_S[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 0.000 2141.670 4.000 ;
    END
  END dyn1_dataIn_S[22]
  PIN dyn1_dataIn_S[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.390 2496.000 2463.670 2500.000 ;
    END
  END dyn1_dataIn_S[23]
  PIN dyn1_dataIn_S[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 2496.000 573.530 2500.000 ;
    END
  END dyn1_dataIn_S[24]
  PIN dyn1_dataIn_S[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 2496.000 393.210 2500.000 ;
    END
  END dyn1_dataIn_S[25]
  PIN dyn1_dataIn_S[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2091.040 4.000 2091.640 ;
    END
  END dyn1_dataIn_S[26]
  PIN dyn1_dataIn_S[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 2496.000 1079.070 2500.000 ;
    END
  END dyn1_dataIn_S[27]
  PIN dyn1_dataIn_S[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 2496.000 1468.690 2500.000 ;
    END
  END dyn1_dataIn_S[28]
  PIN dyn1_dataIn_S[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END dyn1_dataIn_S[29]
  PIN dyn1_dataIn_S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.290 2496.000 1803.570 2500.000 ;
    END
  END dyn1_dataIn_S[2]
  PIN dyn1_dataIn_S[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1329.440 2500.000 1330.040 ;
    END
  END dyn1_dataIn_S[30]
  PIN dyn1_dataIn_S[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 2496.000 145.270 2500.000 ;
    END
  END dyn1_dataIn_S[31]
  PIN dyn1_dataIn_S[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 2496.000 80.870 2500.000 ;
    END
  END dyn1_dataIn_S[32]
  PIN dyn1_dataIn_S[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.110 0.000 2386.390 4.000 ;
    END
  END dyn1_dataIn_S[33]
  PIN dyn1_dataIn_S[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END dyn1_dataIn_S[34]
  PIN dyn1_dataIn_S[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2288.240 4.000 2288.840 ;
    END
  END dyn1_dataIn_S[35]
  PIN dyn1_dataIn_S[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END dyn1_dataIn_S[36]
  PIN dyn1_dataIn_S[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.270 2496.000 2154.550 2500.000 ;
    END
  END dyn1_dataIn_S[37]
  PIN dyn1_dataIn_S[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END dyn1_dataIn_S[38]
  PIN dyn1_dataIn_S[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 2496.000 451.170 2500.000 ;
    END
  END dyn1_dataIn_S[39]
  PIN dyn1_dataIn_S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2060.440 4.000 2061.040 ;
    END
  END dyn1_dataIn_S[3]
  PIN dyn1_dataIn_S[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END dyn1_dataIn_S[40]
  PIN dyn1_dataIn_S[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 2496.000 1529.870 2500.000 ;
    END
  END dyn1_dataIn_S[41]
  PIN dyn1_dataIn_S[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END dyn1_dataIn_S[42]
  PIN dyn1_dataIn_S[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1557.240 4.000 1557.840 ;
    END
  END dyn1_dataIn_S[43]
  PIN dyn1_dataIn_S[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END dyn1_dataIn_S[44]
  PIN dyn1_dataIn_S[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.930 2496.000 2486.210 2500.000 ;
    END
  END dyn1_dataIn_S[45]
  PIN dyn1_dataIn_S[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1057.440 2500.000 1058.040 ;
    END
  END dyn1_dataIn_S[46]
  PIN dyn1_dataIn_S[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END dyn1_dataIn_S[47]
  PIN dyn1_dataIn_S[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 724.240 2500.000 724.840 ;
    END
  END dyn1_dataIn_S[48]
  PIN dyn1_dataIn_S[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 2496.000 563.870 2500.000 ;
    END
  END dyn1_dataIn_S[49]
  PIN dyn1_dataIn_S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END dyn1_dataIn_S[4]
  PIN dyn1_dataIn_S[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 2496.000 608.950 2500.000 ;
    END
  END dyn1_dataIn_S[50]
  PIN dyn1_dataIn_S[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2118.240 2500.000 2118.840 ;
    END
  END dyn1_dataIn_S[51]
  PIN dyn1_dataIn_S[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1125.440 2500.000 1126.040 ;
    END
  END dyn1_dataIn_S[52]
  PIN dyn1_dataIn_S[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 95.240 2500.000 95.840 ;
    END
  END dyn1_dataIn_S[53]
  PIN dyn1_dataIn_S[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1632.040 2500.000 1632.640 ;
    END
  END dyn1_dataIn_S[54]
  PIN dyn1_dataIn_S[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 907.840 2500.000 908.440 ;
    END
  END dyn1_dataIn_S[55]
  PIN dyn1_dataIn_S[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2421.530 0.000 2421.810 4.000 ;
    END
  END dyn1_dataIn_S[56]
  PIN dyn1_dataIn_S[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 0.000 2247.930 4.000 ;
    END
  END dyn1_dataIn_S[57]
  PIN dyn1_dataIn_S[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 329.840 2500.000 330.440 ;
    END
  END dyn1_dataIn_S[58]
  PIN dyn1_dataIn_S[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1577.640 2500.000 1578.240 ;
    END
  END dyn1_dataIn_S[59]
  PIN dyn1_dataIn_S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END dyn1_dataIn_S[5]
  PIN dyn1_dataIn_S[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END dyn1_dataIn_S[60]
  PIN dyn1_dataIn_S[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2036.640 4.000 2037.240 ;
    END
  END dyn1_dataIn_S[61]
  PIN dyn1_dataIn_S[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 697.040 2500.000 697.640 ;
    END
  END dyn1_dataIn_S[62]
  PIN dyn1_dataIn_S[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END dyn1_dataIn_S[63]
  PIN dyn1_dataIn_S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2312.040 4.000 2312.640 ;
    END
  END dyn1_dataIn_S[6]
  PIN dyn1_dataIn_S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2101.240 4.000 2101.840 ;
    END
  END dyn1_dataIn_S[7]
  PIN dyn1_dataIn_S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 2496.000 1871.190 2500.000 ;
    END
  END dyn1_dataIn_S[8]
  PIN dyn1_dataIn_S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1900.640 2500.000 1901.240 ;
    END
  END dyn1_dataIn_S[9]
  PIN dyn1_dataIn_W[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.170 0.000 1977.450 4.000 ;
    END
  END dyn1_dataIn_W[0]
  PIN dyn1_dataIn_W[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END dyn1_dataIn_W[10]
  PIN dyn1_dataIn_W[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END dyn1_dataIn_W[11]
  PIN dyn1_dataIn_W[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 2496.000 1980.670 2500.000 ;
    END
  END dyn1_dataIn_W[12]
  PIN dyn1_dataIn_W[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END dyn1_dataIn_W[13]
  PIN dyn1_dataIn_W[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1761.240 2500.000 1761.840 ;
    END
  END dyn1_dataIn_W[14]
  PIN dyn1_dataIn_W[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END dyn1_dataIn_W[15]
  PIN dyn1_dataIn_W[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2465.040 4.000 2465.640 ;
    END
  END dyn1_dataIn_W[16]
  PIN dyn1_dataIn_W[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 2496.000 827.910 2500.000 ;
    END
  END dyn1_dataIn_W[17]
  PIN dyn1_dataIn_W[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END dyn1_dataIn_W[18]
  PIN dyn1_dataIn_W[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2318.840 4.000 2319.440 ;
    END
  END dyn1_dataIn_W[19]
  PIN dyn1_dataIn_W[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END dyn1_dataIn_W[1]
  PIN dyn1_dataIn_W[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 2496.000 1056.530 2500.000 ;
    END
  END dyn1_dataIn_W[20]
  PIN dyn1_dataIn_W[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END dyn1_dataIn_W[21]
  PIN dyn1_dataIn_W[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 2496.000 769.950 2500.000 ;
    END
  END dyn1_dataIn_W[22]
  PIN dyn1_dataIn_W[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2254.240 4.000 2254.840 ;
    END
  END dyn1_dataIn_W[23]
  PIN dyn1_dataIn_W[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.910 0.000 2032.190 4.000 ;
    END
  END dyn1_dataIn_W[24]
  PIN dyn1_dataIn_W[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1020.040 2500.000 1020.640 ;
    END
  END dyn1_dataIn_W[25]
  PIN dyn1_dataIn_W[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 2496.000 670.130 2500.000 ;
    END
  END dyn1_dataIn_W[26]
  PIN dyn1_dataIn_W[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 0.000 1401.070 4.000 ;
    END
  END dyn1_dataIn_W[27]
  PIN dyn1_dataIn_W[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 2496.000 998.570 2500.000 ;
    END
  END dyn1_dataIn_W[28]
  PIN dyn1_dataIn_W[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END dyn1_dataIn_W[29]
  PIN dyn1_dataIn_W[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1781.640 2500.000 1782.240 ;
    END
  END dyn1_dataIn_W[2]
  PIN dyn1_dataIn_W[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END dyn1_dataIn_W[30]
  PIN dyn1_dataIn_W[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 2496.000 1674.770 2500.000 ;
    END
  END dyn1_dataIn_W[31]
  PIN dyn1_dataIn_W[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.040 4.000 1632.640 ;
    END
  END dyn1_dataIn_W[32]
  PIN dyn1_dataIn_W[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 0.000 2112.690 4.000 ;
    END
  END dyn1_dataIn_W[33]
  PIN dyn1_dataIn_W[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1390.640 2500.000 1391.240 ;
    END
  END dyn1_dataIn_W[34]
  PIN dyn1_dataIn_W[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END dyn1_dataIn_W[35]
  PIN dyn1_dataIn_W[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END dyn1_dataIn_W[36]
  PIN dyn1_dataIn_W[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 2496.000 212.890 2500.000 ;
    END
  END dyn1_dataIn_W[37]
  PIN dyn1_dataIn_W[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1703.440 2500.000 1704.040 ;
    END
  END dyn1_dataIn_W[38]
  PIN dyn1_dataIn_W[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2067.240 4.000 2067.840 ;
    END
  END dyn1_dataIn_W[39]
  PIN dyn1_dataIn_W[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 2496.000 1043.650 2500.000 ;
    END
  END dyn1_dataIn_W[3]
  PIN dyn1_dataIn_W[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END dyn1_dataIn_W[40]
  PIN dyn1_dataIn_W[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.950 0.000 2457.230 4.000 ;
    END
  END dyn1_dataIn_W[41]
  PIN dyn1_dataIn_W[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 506.640 2500.000 507.240 ;
    END
  END dyn1_dataIn_W[42]
  PIN dyn1_dataIn_W[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 666.440 2500.000 667.040 ;
    END
  END dyn1_dataIn_W[43]
  PIN dyn1_dataIn_W[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1904.040 4.000 1904.640 ;
    END
  END dyn1_dataIn_W[44]
  PIN dyn1_dataIn_W[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2465.040 2500.000 2465.640 ;
    END
  END dyn1_dataIn_W[45]
  PIN dyn1_dataIn_W[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END dyn1_dataIn_W[46]
  PIN dyn1_dataIn_W[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 2496.000 528.450 2500.000 ;
    END
  END dyn1_dataIn_W[47]
  PIN dyn1_dataIn_W[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1479.040 2500.000 1479.640 ;
    END
  END dyn1_dataIn_W[48]
  PIN dyn1_dataIn_W[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 2496.000 583.190 2500.000 ;
    END
  END dyn1_dataIn_W[49]
  PIN dyn1_dataIn_W[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 2496.000 853.670 2500.000 ;
    END
  END dyn1_dataIn_W[4]
  PIN dyn1_dataIn_W[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END dyn1_dataIn_W[50]
  PIN dyn1_dataIn_W[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.970 2496.000 2267.250 2500.000 ;
    END
  END dyn1_dataIn_W[51]
  PIN dyn1_dataIn_W[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1343.040 2500.000 1343.640 ;
    END
  END dyn1_dataIn_W[52]
  PIN dyn1_dataIn_W[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1509.640 2500.000 1510.240 ;
    END
  END dyn1_dataIn_W[53]
  PIN dyn1_dataIn_W[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END dyn1_dataIn_W[54]
  PIN dyn1_dataIn_W[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END dyn1_dataIn_W[55]
  PIN dyn1_dataIn_W[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2444.640 2500.000 2445.240 ;
    END
  END dyn1_dataIn_W[56]
  PIN dyn1_dataIn_W[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 2496.000 1748.830 2500.000 ;
    END
  END dyn1_dataIn_W[57]
  PIN dyn1_dataIn_W[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 248.240 2500.000 248.840 ;
    END
  END dyn1_dataIn_W[58]
  PIN dyn1_dataIn_W[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 992.840 2500.000 993.440 ;
    END
  END dyn1_dataIn_W[59]
  PIN dyn1_dataIn_W[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END dyn1_dataIn_W[5]
  PIN dyn1_dataIn_W[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2029.840 2500.000 2030.440 ;
    END
  END dyn1_dataIn_W[60]
  PIN dyn1_dataIn_W[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END dyn1_dataIn_W[61]
  PIN dyn1_dataIn_W[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END dyn1_dataIn_W[62]
  PIN dyn1_dataIn_W[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 2496.000 1855.090 2500.000 ;
    END
  END dyn1_dataIn_W[63]
  PIN dyn1_dataIn_W[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END dyn1_dataIn_W[6]
  PIN dyn1_dataIn_W[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2104.640 2500.000 2105.240 ;
    END
  END dyn1_dataIn_W[7]
  PIN dyn1_dataIn_W[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 2496.000 641.150 2500.000 ;
    END
  END dyn1_dataIn_W[8]
  PIN dyn1_dataIn_W[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1060.840 2500.000 1061.440 ;
    END
  END dyn1_dataIn_W[9]
  PIN dyn1_validIn_E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.570 2496.000 2041.850 2500.000 ;
    END
  END dyn1_validIn_E
  PIN dyn1_validIn_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END dyn1_validIn_N
  PIN dyn1_validIn_S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.290 0.000 1964.570 4.000 ;
    END
  END dyn1_validIn_S
  PIN dyn1_validIn_W
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2261.040 2500.000 2261.640 ;
    END
  END dyn1_validIn_W
  PIN dyn1_yummyOut_E
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1152.640 2500.000 1153.240 ;
    END
  END dyn1_yummyOut_E
  PIN dyn1_yummyOut_N
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END dyn1_yummyOut_N
  PIN dyn1_yummyOut_S
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 2496.000 1887.290 2500.000 ;
    END
  END dyn1_yummyOut_S
  PIN dyn1_yummyOut_W
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END dyn1_yummyOut_W
  PIN dyn2_dEo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 2496.000 1059.750 2500.000 ;
    END
  END dyn2_dEo[0]
  PIN dyn2_dEo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 0.000 1684.430 4.000 ;
    END
  END dyn2_dEo[10]
  PIN dyn2_dEo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1414.440 2500.000 1415.040 ;
    END
  END dyn2_dEo[11]
  PIN dyn2_dEo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1533.440 4.000 1534.040 ;
    END
  END dyn2_dEo[12]
  PIN dyn2_dEo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2499.040 4.000 2499.640 ;
    END
  END dyn2_dEo[13]
  PIN dyn2_dEo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 2496.000 209.670 2500.000 ;
    END
  END dyn2_dEo[14]
  PIN dyn2_dEo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 2496.000 1520.210 2500.000 ;
    END
  END dyn2_dEo[15]
  PIN dyn2_dEo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 2496.000 1929.150 2500.000 ;
    END
  END dyn2_dEo[16]
  PIN dyn2_dEo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 2496.000 657.250 2500.000 ;
    END
  END dyn2_dEo[17]
  PIN dyn2_dEo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 2496.000 689.450 2500.000 ;
    END
  END dyn2_dEo[18]
  PIN dyn2_dEo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END dyn2_dEo[19]
  PIN dyn2_dEo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END dyn2_dEo[1]
  PIN dyn2_dEo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END dyn2_dEo[20]
  PIN dyn2_dEo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 0.000 1240.070 4.000 ;
    END
  END dyn2_dEo[21]
  PIN dyn2_dEo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END dyn2_dEo[22]
  PIN dyn2_dEo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END dyn2_dEo[23]
  PIN dyn2_dEo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 890.840 2500.000 891.440 ;
    END
  END dyn2_dEo[24]
  PIN dyn2_dEo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 4.000 ;
    END
  END dyn2_dEo[25]
  PIN dyn2_dEo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END dyn2_dEo[26]
  PIN dyn2_dEo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2475.240 2500.000 2475.840 ;
    END
  END dyn2_dEo[27]
  PIN dyn2_dEo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.610 2496.000 2466.890 2500.000 ;
    END
  END dyn2_dEo[28]
  PIN dyn2_dEo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END dyn2_dEo[29]
  PIN dyn2_dEo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END dyn2_dEo[2]
  PIN dyn2_dEo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END dyn2_dEo[30]
  PIN dyn2_dEo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.550 0.000 2231.830 4.000 ;
    END
  END dyn2_dEo[31]
  PIN dyn2_dEo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 2496.000 354.570 2500.000 ;
    END
  END dyn2_dEo[32]
  PIN dyn2_dEo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.330 2496.000 2067.610 2500.000 ;
    END
  END dyn2_dEo[33]
  PIN dyn2_dEo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END dyn2_dEo[34]
  PIN dyn2_dEo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 448.840 2500.000 449.440 ;
    END
  END dyn2_dEo[35]
  PIN dyn2_dEo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 2496.000 306.270 2500.000 ;
    END
  END dyn2_dEo[36]
  PIN dyn2_dEo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 2496.000 686.230 2500.000 ;
    END
  END dyn2_dEo[37]
  PIN dyn2_dEo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.230 0.000 2373.510 4.000 ;
    END
  END dyn2_dEo[38]
  PIN dyn2_dEo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2220.240 2500.000 2220.840 ;
    END
  END dyn2_dEo[39]
  PIN dyn2_dEo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END dyn2_dEo[3]
  PIN dyn2_dEo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END dyn2_dEo[40]
  PIN dyn2_dEo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 2496.000 618.610 2500.000 ;
    END
  END dyn2_dEo[41]
  PIN dyn2_dEo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END dyn2_dEo[42]
  PIN dyn2_dEo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END dyn2_dEo[43]
  PIN dyn2_dEo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1380.440 2500.000 1381.040 ;
    END
  END dyn2_dEo[44]
  PIN dyn2_dEo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 557.640 2500.000 558.240 ;
    END
  END dyn2_dEo[45]
  PIN dyn2_dEo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2169.240 4.000 2169.840 ;
    END
  END dyn2_dEo[46]
  PIN dyn2_dEo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2012.840 4.000 2013.440 ;
    END
  END dyn2_dEo[47]
  PIN dyn2_dEo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END dyn2_dEo[48]
  PIN dyn2_dEo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END dyn2_dEo[49]
  PIN dyn2_dEo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1230.840 2500.000 1231.440 ;
    END
  END dyn2_dEo[4]
  PIN dyn2_dEo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.310 2496.000 2096.590 2500.000 ;
    END
  END dyn2_dEo[50]
  PIN dyn2_dEo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END dyn2_dEo[51]
  PIN dyn2_dEo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 4.000 ;
    END
  END dyn2_dEo[52]
  PIN dyn2_dEo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END dyn2_dEo[53]
  PIN dyn2_dEo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 4.000 ;
    END
  END dyn2_dEo[54]
  PIN dyn2_dEo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 2496.000 2183.530 2500.000 ;
    END
  END dyn2_dEo[55]
  PIN dyn2_dEo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END dyn2_dEo[56]
  PIN dyn2_dEo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 0.000 1027.550 4.000 ;
    END
  END dyn2_dEo[57]
  PIN dyn2_dEo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1431.440 2500.000 1432.040 ;
    END
  END dyn2_dEo[58]
  PIN dyn2_dEo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1802.040 2500.000 1802.640 ;
    END
  END dyn2_dEo[59]
  PIN dyn2_dEo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 4.000 ;
    END
  END dyn2_dEo[5]
  PIN dyn2_dEo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END dyn2_dEo[60]
  PIN dyn2_dEo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 391.040 2500.000 391.640 ;
    END
  END dyn2_dEo[61]
  PIN dyn2_dEo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 197.240 2500.000 197.840 ;
    END
  END dyn2_dEo[62]
  PIN dyn2_dEo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 316.240 2500.000 316.840 ;
    END
  END dyn2_dEo[63]
  PIN dyn2_dEo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1176.440 2500.000 1177.040 ;
    END
  END dyn2_dEo[6]
  PIN dyn2_dEo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2305.240 2500.000 2305.840 ;
    END
  END dyn2_dEo[7]
  PIN dyn2_dEo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2305.610 2496.000 2305.890 2500.000 ;
    END
  END dyn2_dEo[8]
  PIN dyn2_dEo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 2496.000 924.510 2500.000 ;
    END
  END dyn2_dEo[9]
  PIN dyn2_dEo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 2496.000 1349.550 2500.000 ;
    END
  END dyn2_dEo_valid
  PIN dyn2_dEo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.710 2496.000 1677.990 2500.000 ;
    END
  END dyn2_dEo_yummy
  PIN dyn2_dNo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 2496.000 676.570 2500.000 ;
    END
  END dyn2_dNo[0]
  PIN dyn2_dNo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END dyn2_dNo[10]
  PIN dyn2_dNo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 2496.000 2431.470 2500.000 ;
    END
  END dyn2_dNo[11]
  PIN dyn2_dNo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1727.240 2500.000 1727.840 ;
    END
  END dyn2_dNo[12]
  PIN dyn2_dNo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END dyn2_dNo[13]
  PIN dyn2_dNo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1995.840 2500.000 1996.440 ;
    END
  END dyn2_dNo[14]
  PIN dyn2_dNo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2274.640 2500.000 2275.240 ;
    END
  END dyn2_dNo[15]
  PIN dyn2_dNo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1999.240 4.000 1999.840 ;
    END
  END dyn2_dNo[16]
  PIN dyn2_dNo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END dyn2_dNo[17]
  PIN dyn2_dNo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 2496.000 332.030 2500.000 ;
    END
  END dyn2_dNo[18]
  PIN dyn2_dNo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 2496.000 1194.990 2500.000 ;
    END
  END dyn2_dNo[19]
  PIN dyn2_dNo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1006.440 4.000 1007.040 ;
    END
  END dyn2_dNo[1]
  PIN dyn2_dNo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.290 2496.000 2286.570 2500.000 ;
    END
  END dyn2_dNo[20]
  PIN dyn2_dNo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.350 2496.000 2360.630 2500.000 ;
    END
  END dyn2_dNo[21]
  PIN dyn2_dNo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1115.240 2500.000 1115.840 ;
    END
  END dyn2_dNo[22]
  PIN dyn2_dNo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 2496.000 879.430 2500.000 ;
    END
  END dyn2_dNo[23]
  PIN dyn2_dNo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END dyn2_dNo[24]
  PIN dyn2_dNo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 190.440 2500.000 191.040 ;
    END
  END dyn2_dNo[25]
  PIN dyn2_dNo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 2496.000 1620.030 2500.000 ;
    END
  END dyn2_dNo[26]
  PIN dyn2_dNo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END dyn2_dNo[27]
  PIN dyn2_dNo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1917.640 2500.000 1918.240 ;
    END
  END dyn2_dNo[28]
  PIN dyn2_dNo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END dyn2_dNo[29]
  PIN dyn2_dNo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END dyn2_dNo[2]
  PIN dyn2_dNo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END dyn2_dNo[30]
  PIN dyn2_dNo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END dyn2_dNo[31]
  PIN dyn2_dNo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END dyn2_dNo[32]
  PIN dyn2_dNo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 2496.000 1845.430 2500.000 ;
    END
  END dyn2_dNo[33]
  PIN dyn2_dNo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END dyn2_dNo[34]
  PIN dyn2_dNo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END dyn2_dNo[35]
  PIN dyn2_dNo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END dyn2_dNo[36]
  PIN dyn2_dNo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2138.640 4.000 2139.240 ;
    END
  END dyn2_dNo[37]
  PIN dyn2_dNo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END dyn2_dNo[38]
  PIN dyn2_dNo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 2496.000 1639.350 2500.000 ;
    END
  END dyn2_dNo[39]
  PIN dyn2_dNo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END dyn2_dNo[3]
  PIN dyn2_dNo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END dyn2_dNo[40]
  PIN dyn2_dNo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END dyn2_dNo[41]
  PIN dyn2_dNo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1992.440 4.000 1993.040 ;
    END
  END dyn2_dNo[42]
  PIN dyn2_dNo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 4.000 ;
    END
  END dyn2_dNo[43]
  PIN dyn2_dNo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2471.840 2500.000 2472.440 ;
    END
  END dyn2_dNo[44]
  PIN dyn2_dNo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 676.640 2500.000 677.240 ;
    END
  END dyn2_dNo[45]
  PIN dyn2_dNo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 0.000 1713.410 4.000 ;
    END
  END dyn2_dNo[46]
  PIN dyn2_dNo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 2496.000 2241.490 2500.000 ;
    END
  END dyn2_dNo[47]
  PIN dyn2_dNo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 91.840 2500.000 92.440 ;
    END
  END dyn2_dNo[48]
  PIN dyn2_dNo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1778.240 4.000 1778.840 ;
    END
  END dyn2_dNo[49]
  PIN dyn2_dNo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END dyn2_dNo[4]
  PIN dyn2_dNo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END dyn2_dNo[50]
  PIN dyn2_dNo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 700.440 2500.000 701.040 ;
    END
  END dyn2_dNo[51]
  PIN dyn2_dNo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 2496.000 1153.130 2500.000 ;
    END
  END dyn2_dNo[52]
  PIN dyn2_dNo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 2496.000 206.450 2500.000 ;
    END
  END dyn2_dNo[53]
  PIN dyn2_dNo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 0.000 1893.730 4.000 ;
    END
  END dyn2_dNo[54]
  PIN dyn2_dNo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2159.040 4.000 2159.640 ;
    END
  END dyn2_dNo[55]
  PIN dyn2_dNo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END dyn2_dNo[56]
  PIN dyn2_dNo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 0.000 1980.670 4.000 ;
    END
  END dyn2_dNo[57]
  PIN dyn2_dNo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END dyn2_dNo[58]
  PIN dyn2_dNo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 479.440 2500.000 480.040 ;
    END
  END dyn2_dNo[59]
  PIN dyn2_dNo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.750 0.000 2264.030 4.000 ;
    END
  END dyn2_dNo[5]
  PIN dyn2_dNo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 2496.000 2103.030 2500.000 ;
    END
  END dyn2_dNo[60]
  PIN dyn2_dNo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.530 2496.000 1938.810 2500.000 ;
    END
  END dyn2_dNo[61]
  PIN dyn2_dNo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END dyn2_dNo[62]
  PIN dyn2_dNo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 2496.000 483.370 2500.000 ;
    END
  END dyn2_dNo[63]
  PIN dyn2_dNo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END dyn2_dNo[6]
  PIN dyn2_dNo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END dyn2_dNo[7]
  PIN dyn2_dNo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 608.640 2500.000 609.240 ;
    END
  END dyn2_dNo[8]
  PIN dyn2_dNo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END dyn2_dNo[9]
  PIN dyn2_dNo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END dyn2_dNo_valid
  PIN dyn2_dNo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 136.040 2500.000 136.640 ;
    END
  END dyn2_dNo_yummy
  PIN dyn2_dSo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 975.840 2500.000 976.440 ;
    END
  END dyn2_dSo[0]
  PIN dyn2_dSo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1764.640 2500.000 1765.240 ;
    END
  END dyn2_dSo[10]
  PIN dyn2_dSo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.350 0.000 1877.630 4.000 ;
    END
  END dyn2_dSo[11]
  PIN dyn2_dSo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1156.040 2500.000 1156.640 ;
    END
  END dyn2_dSo[12]
  PIN dyn2_dSo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 2496.000 728.090 2500.000 ;
    END
  END dyn2_dSo[13]
  PIN dyn2_dSo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 680.040 2500.000 680.640 ;
    END
  END dyn2_dSo[14]
  PIN dyn2_dSo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END dyn2_dSo[15]
  PIN dyn2_dSo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END dyn2_dSo[16]
  PIN dyn2_dSo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 2496.000 1333.450 2500.000 ;
    END
  END dyn2_dSo[17]
  PIN dyn2_dSo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END dyn2_dSo[18]
  PIN dyn2_dSo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1900.640 4.000 1901.240 ;
    END
  END dyn2_dSo[19]
  PIN dyn2_dSo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 4.000 ;
    END
  END dyn2_dSo[1]
  PIN dyn2_dSo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 2496.000 918.070 2500.000 ;
    END
  END dyn2_dSo[20]
  PIN dyn2_dSo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 0.000 1124.150 4.000 ;
    END
  END dyn2_dSo[21]
  PIN dyn2_dSo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2091.040 2500.000 2091.640 ;
    END
  END dyn2_dSo[22]
  PIN dyn2_dSo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END dyn2_dSo[23]
  PIN dyn2_dSo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END dyn2_dSo[24]
  PIN dyn2_dSo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2410.640 4.000 2411.240 ;
    END
  END dyn2_dSo[25]
  PIN dyn2_dSo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END dyn2_dSo[26]
  PIN dyn2_dSo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 2496.000 489.810 2500.000 ;
    END
  END dyn2_dSo[27]
  PIN dyn2_dSo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 2496.000 612.170 2500.000 ;
    END
  END dyn2_dSo[28]
  PIN dyn2_dSo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END dyn2_dSo[29]
  PIN dyn2_dSo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1876.840 4.000 1877.440 ;
    END
  END dyn2_dSo[2]
  PIN dyn2_dSo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2451.440 4.000 2452.040 ;
    END
  END dyn2_dSo[30]
  PIN dyn2_dSo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.510 0.000 2128.790 4.000 ;
    END
  END dyn2_dSo[31]
  PIN dyn2_dSo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 377.440 2500.000 378.040 ;
    END
  END dyn2_dSo[32]
  PIN dyn2_dSo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 0.000 1903.390 4.000 ;
    END
  END dyn2_dSo[33]
  PIN dyn2_dSo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.210 0.000 2402.490 4.000 ;
    END
  END dyn2_dSo[34]
  PIN dyn2_dSo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 2496.000 589.630 2500.000 ;
    END
  END dyn2_dSo[35]
  PIN dyn2_dSo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END dyn2_dSo[36]
  PIN dyn2_dSo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 2496.000 1172.450 2500.000 ;
    END
  END dyn2_dSo[37]
  PIN dyn2_dSo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 384.240 2500.000 384.840 ;
    END
  END dyn2_dSo[38]
  PIN dyn2_dSo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1625.240 2500.000 1625.840 ;
    END
  END dyn2_dSo[39]
  PIN dyn2_dSo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 272.040 2500.000 272.640 ;
    END
  END dyn2_dSo[3]
  PIN dyn2_dSo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2172.640 2500.000 2173.240 ;
    END
  END dyn2_dSo[40]
  PIN dyn2_dSo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.840 4.000 1486.440 ;
    END
  END dyn2_dSo[41]
  PIN dyn2_dSo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END dyn2_dSo[42]
  PIN dyn2_dSo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1434.840 2500.000 1435.440 ;
    END
  END dyn2_dSo[43]
  PIN dyn2_dSo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 2496.000 6.810 2500.000 ;
    END
  END dyn2_dSo[44]
  PIN dyn2_dSo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 0.000 1365.650 4.000 ;
    END
  END dyn2_dSo[45]
  PIN dyn2_dSo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 2496.000 1494.450 2500.000 ;
    END
  END dyn2_dSo[46]
  PIN dyn2_dSo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1720.440 4.000 1721.040 ;
    END
  END dyn2_dSo[47]
  PIN dyn2_dSo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END dyn2_dSo[48]
  PIN dyn2_dSo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END dyn2_dSo[49]
  PIN dyn2_dSo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1492.640 2500.000 1493.240 ;
    END
  END dyn2_dSo[4]
  PIN dyn2_dSo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 2496.000 995.350 2500.000 ;
    END
  END dyn2_dSo[50]
  PIN dyn2_dSo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END dyn2_dSo[51]
  PIN dyn2_dSo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1761.240 4.000 1761.840 ;
    END
  END dyn2_dSo[52]
  PIN dyn2_dSo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 2496.000 493.030 2500.000 ;
    END
  END dyn2_dSo[53]
  PIN dyn2_dSo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 914.640 2500.000 915.240 ;
    END
  END dyn2_dSo[54]
  PIN dyn2_dSo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 0.000 1288.370 4.000 ;
    END
  END dyn2_dSo[55]
  PIN dyn2_dSo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 149.640 2500.000 150.240 ;
    END
  END dyn2_dSo[56]
  PIN dyn2_dSo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END dyn2_dSo[57]
  PIN dyn2_dSo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END dyn2_dSo[58]
  PIN dyn2_dSo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.840 4.000 1418.440 ;
    END
  END dyn2_dSo[59]
  PIN dyn2_dSo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END dyn2_dSo[5]
  PIN dyn2_dSo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.510 2496.000 1967.790 2500.000 ;
    END
  END dyn2_dSo[60]
  PIN dyn2_dSo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END dyn2_dSo[61]
  PIN dyn2_dSo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 812.640 2500.000 813.240 ;
    END
  END dyn2_dSo[62]
  PIN dyn2_dSo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1693.240 2500.000 1693.840 ;
    END
  END dyn2_dSo[63]
  PIN dyn2_dSo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END dyn2_dSo[6]
  PIN dyn2_dSo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2033.240 2500.000 2033.840 ;
    END
  END dyn2_dSo[7]
  PIN dyn2_dSo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2400.440 2500.000 2401.040 ;
    END
  END dyn2_dSo[8]
  PIN dyn2_dSo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2009.440 4.000 2010.040 ;
    END
  END dyn2_dSo[9]
  PIN dyn2_dSo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END dyn2_dSo_valid
  PIN dyn2_dSo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 2496.000 16.470 2500.000 ;
    END
  END dyn2_dSo_yummy
  PIN dyn2_dWo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END dyn2_dWo[0]
  PIN dyn2_dWo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 2496.000 2293.010 2500.000 ;
    END
  END dyn2_dWo[10]
  PIN dyn2_dWo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END dyn2_dWo[11]
  PIN dyn2_dWo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 2496.000 51.890 2500.000 ;
    END
  END dyn2_dWo[12]
  PIN dyn2_dWo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 2496.000 1632.910 2500.000 ;
    END
  END dyn2_dWo[13]
  PIN dyn2_dWo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END dyn2_dWo[14]
  PIN dyn2_dWo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1377.040 2500.000 1377.640 ;
    END
  END dyn2_dWo[15]
  PIN dyn2_dWo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1026.840 2500.000 1027.440 ;
    END
  END dyn2_dWo[16]
  PIN dyn2_dWo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 170.040 2500.000 170.640 ;
    END
  END dyn2_dWo[17]
  PIN dyn2_dWo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2036.640 2500.000 2037.240 ;
    END
  END dyn2_dWo[18]
  PIN dyn2_dWo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END dyn2_dWo[19]
  PIN dyn2_dWo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END dyn2_dWo[1]
  PIN dyn2_dWo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END dyn2_dWo[20]
  PIN dyn2_dWo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END dyn2_dWo[21]
  PIN dyn2_dWo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END dyn2_dWo[22]
  PIN dyn2_dWo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END dyn2_dWo[23]
  PIN dyn2_dWo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END dyn2_dWo[24]
  PIN dyn2_dWo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.470 0.000 2025.750 4.000 ;
    END
  END dyn2_dWo[25]
  PIN dyn2_dWo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.110 2496.000 2386.390 2500.000 ;
    END
  END dyn2_dWo[26]
  PIN dyn2_dWo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END dyn2_dWo[27]
  PIN dyn2_dWo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 0.000 1983.890 4.000 ;
    END
  END dyn2_dWo[28]
  PIN dyn2_dWo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 74.840 2500.000 75.440 ;
    END
  END dyn2_dWo[29]
  PIN dyn2_dWo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END dyn2_dWo[2]
  PIN dyn2_dWo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END dyn2_dWo[30]
  PIN dyn2_dWo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 2496.000 1661.890 2500.000 ;
    END
  END dyn2_dWo[31]
  PIN dyn2_dWo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END dyn2_dWo[32]
  PIN dyn2_dWo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END dyn2_dWo[33]
  PIN dyn2_dWo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END dyn2_dWo[34]
  PIN dyn2_dWo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 2496.000 1082.290 2500.000 ;
    END
  END dyn2_dWo[35]
  PIN dyn2_dWo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 2496.000 660.470 2500.000 ;
    END
  END dyn2_dWo[36]
  PIN dyn2_dWo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1802.040 4.000 1802.640 ;
    END
  END dyn2_dWo[37]
  PIN dyn2_dWo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END dyn2_dWo[38]
  PIN dyn2_dWo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 2496.000 1207.870 2500.000 ;
    END
  END dyn2_dWo[39]
  PIN dyn2_dWo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END dyn2_dWo[3]
  PIN dyn2_dWo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END dyn2_dWo[40]
  PIN dyn2_dWo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END dyn2_dWo[41]
  PIN dyn2_dWo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.840 4.000 1282.440 ;
    END
  END dyn2_dWo[42]
  PIN dyn2_dWo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 2496.000 586.410 2500.000 ;
    END
  END dyn2_dWo[43]
  PIN dyn2_dWo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 2496.000 1880.850 2500.000 ;
    END
  END dyn2_dWo[44]
  PIN dyn2_dWo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END dyn2_dWo[45]
  PIN dyn2_dWo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 2496.000 319.150 2500.000 ;
    END
  END dyn2_dWo[46]
  PIN dyn2_dWo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 187.040 2500.000 187.640 ;
    END
  END dyn2_dWo[47]
  PIN dyn2_dWo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.750 2496.000 2425.030 2500.000 ;
    END
  END dyn2_dWo[48]
  PIN dyn2_dWo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 2496.000 1417.170 2500.000 ;
    END
  END dyn2_dWo[49]
  PIN dyn2_dWo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END dyn2_dWo[4]
  PIN dyn2_dWo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1560.640 4.000 1561.240 ;
    END
  END dyn2_dWo[50]
  PIN dyn2_dWo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 2496.000 866.550 2500.000 ;
    END
  END dyn2_dWo[51]
  PIN dyn2_dWo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END dyn2_dWo[52]
  PIN dyn2_dWo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 2496.000 1169.230 2500.000 ;
    END
  END dyn2_dWo[53]
  PIN dyn2_dWo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1203.640 2500.000 1204.240 ;
    END
  END dyn2_dWo[54]
  PIN dyn2_dWo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1543.640 2500.000 1544.240 ;
    END
  END dyn2_dWo[55]
  PIN dyn2_dWo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END dyn2_dWo[56]
  PIN dyn2_dWo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 2496.000 1050.090 2500.000 ;
    END
  END dyn2_dWo[57]
  PIN dyn2_dWo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2417.440 4.000 2418.040 ;
    END
  END dyn2_dWo[58]
  PIN dyn2_dWo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 2496.000 1433.270 2500.000 ;
    END
  END dyn2_dWo[59]
  PIN dyn2_dWo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END dyn2_dWo[5]
  PIN dyn2_dWo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 2496.000 228.990 2500.000 ;
    END
  END dyn2_dWo[60]
  PIN dyn2_dWo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 2496.000 663.690 2500.000 ;
    END
  END dyn2_dWo[61]
  PIN dyn2_dWo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 595.040 2500.000 595.640 ;
    END
  END dyn2_dWo[62]
  PIN dyn2_dWo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END dyn2_dWo[63]
  PIN dyn2_dWo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END dyn2_dWo[6]
  PIN dyn2_dWo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 2496.000 1355.990 2500.000 ;
    END
  END dyn2_dWo[7]
  PIN dyn2_dWo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END dyn2_dWo[8]
  PIN dyn2_dWo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 2496.000 438.290 2500.000 ;
    END
  END dyn2_dWo[9]
  PIN dyn2_dWo_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END dyn2_dWo_valid
  PIN dyn2_dWo_yummy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END dyn2_dWo_yummy
  PIN dyn2_dataIn_E[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END dyn2_dataIn_E[0]
  PIN dyn2_dataIn_E[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 343.440 2500.000 344.040 ;
    END
  END dyn2_dataIn_E[10]
  PIN dyn2_dataIn_E[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 2496.000 1510.550 2500.000 ;
    END
  END dyn2_dataIn_E[11]
  PIN dyn2_dataIn_E[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 2496.000 1739.170 2500.000 ;
    END
  END dyn2_dataIn_E[12]
  PIN dyn2_dataIn_E[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END dyn2_dataIn_E[13]
  PIN dyn2_dataIn_E[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 146.240 2500.000 146.840 ;
    END
  END dyn2_dataIn_E[14]
  PIN dyn2_dataIn_E[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END dyn2_dataIn_E[15]
  PIN dyn2_dataIn_E[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END dyn2_dataIn_E[16]
  PIN dyn2_dataIn_E[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2040.040 2500.000 2040.640 ;
    END
  END dyn2_dataIn_E[17]
  PIN dyn2_dataIn_E[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1944.840 4.000 1945.440 ;
    END
  END dyn2_dataIn_E[18]
  PIN dyn2_dataIn_E[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2488.840 2500.000 2489.440 ;
    END
  END dyn2_dataIn_E[19]
  PIN dyn2_dataIn_E[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 2496.000 32.570 2500.000 ;
    END
  END dyn2_dataIn_E[1]
  PIN dyn2_dataIn_E[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 159.840 2500.000 160.440 ;
    END
  END dyn2_dataIn_E[20]
  PIN dyn2_dataIn_E[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END dyn2_dataIn_E[21]
  PIN dyn2_dataIn_E[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 2496.000 1404.290 2500.000 ;
    END
  END dyn2_dataIn_E[22]
  PIN dyn2_dataIn_E[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2019.640 4.000 2020.240 ;
    END
  END dyn2_dataIn_E[23]
  PIN dyn2_dataIn_E[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1621.840 2500.000 1622.440 ;
    END
  END dyn2_dataIn_E[24]
  PIN dyn2_dataIn_E[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.230 2496.000 2373.510 2500.000 ;
    END
  END dyn2_dataIn_E[25]
  PIN dyn2_dataIn_E[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2240.640 4.000 2241.240 ;
    END
  END dyn2_dataIn_E[26]
  PIN dyn2_dataIn_E[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1169.640 2500.000 1170.240 ;
    END
  END dyn2_dataIn_E[27]
  PIN dyn2_dataIn_E[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END dyn2_dataIn_E[28]
  PIN dyn2_dataIn_E[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.170 0.000 2299.450 4.000 ;
    END
  END dyn2_dataIn_E[29]
  PIN dyn2_dataIn_E[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 2496.000 2077.270 2500.000 ;
    END
  END dyn2_dataIn_E[2]
  PIN dyn2_dataIn_E[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2169.240 2500.000 2169.840 ;
    END
  END dyn2_dataIn_E[30]
  PIN dyn2_dataIn_E[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 129.240 2500.000 129.840 ;
    END
  END dyn2_dataIn_E[31]
  PIN dyn2_dataIn_E[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 516.840 2500.000 517.440 ;
    END
  END dyn2_dataIn_E[32]
  PIN dyn2_dataIn_E[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 727.640 2500.000 728.240 ;
    END
  END dyn2_dataIn_E[33]
  PIN dyn2_dataIn_E[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.690 0.000 2028.970 4.000 ;
    END
  END dyn2_dataIn_E[34]
  PIN dyn2_dataIn_E[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1832.640 2500.000 1833.240 ;
    END
  END dyn2_dataIn_E[35]
  PIN dyn2_dataIn_E[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 2496.000 1359.210 2500.000 ;
    END
  END dyn2_dataIn_E[36]
  PIN dyn2_dataIn_E[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END dyn2_dataIn_E[37]
  PIN dyn2_dataIn_E[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1921.040 4.000 1921.640 ;
    END
  END dyn2_dataIn_E[38]
  PIN dyn2_dataIn_E[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 782.040 2500.000 782.640 ;
    END
  END dyn2_dataIn_E[39]
  PIN dyn2_dataIn_E[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 0.000 2293.010 4.000 ;
    END
  END dyn2_dataIn_E[3]
  PIN dyn2_dataIn_E[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1292.040 2500.000 1292.640 ;
    END
  END dyn2_dataIn_E[40]
  PIN dyn2_dataIn_E[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1006.440 2500.000 1007.040 ;
    END
  END dyn2_dataIn_E[41]
  PIN dyn2_dataIn_E[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1122.040 2500.000 1122.640 ;
    END
  END dyn2_dataIn_E[42]
  PIN dyn2_dataIn_E[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1149.240 4.000 1149.840 ;
    END
  END dyn2_dataIn_E[43]
  PIN dyn2_dataIn_E[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 2496.000 129.170 2500.000 ;
    END
  END dyn2_dataIn_E[44]
  PIN dyn2_dataIn_E[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 2496.000 1256.170 2500.000 ;
    END
  END dyn2_dataIn_E[45]
  PIN dyn2_dataIn_E[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1186.640 2500.000 1187.240 ;
    END
  END dyn2_dataIn_E[46]
  PIN dyn2_dataIn_E[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END dyn2_dataIn_E[47]
  PIN dyn2_dataIn_E[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.670 2496.000 2057.950 2500.000 ;
    END
  END dyn2_dataIn_E[48]
  PIN dyn2_dataIn_E[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 2496.000 290.170 2500.000 ;
    END
  END dyn2_dataIn_E[49]
  PIN dyn2_dataIn_E[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2363.040 2500.000 2363.640 ;
    END
  END dyn2_dataIn_E[4]
  PIN dyn2_dataIn_E[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1737.440 2500.000 1738.040 ;
    END
  END dyn2_dataIn_E[50]
  PIN dyn2_dataIn_E[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END dyn2_dataIn_E[51]
  PIN dyn2_dataIn_E[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END dyn2_dataIn_E[52]
  PIN dyn2_dataIn_E[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2247.440 2500.000 2248.040 ;
    END
  END dyn2_dataIn_E[53]
  PIN dyn2_dataIn_E[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.240 4.000 1608.840 ;
    END
  END dyn2_dataIn_E[54]
  PIN dyn2_dataIn_E[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.710 0.000 2482.990 4.000 ;
    END
  END dyn2_dataIn_E[55]
  PIN dyn2_dataIn_E[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END dyn2_dataIn_E[56]
  PIN dyn2_dataIn_E[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END dyn2_dataIn_E[57]
  PIN dyn2_dataIn_E[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 2496.000 579.970 2500.000 ;
    END
  END dyn2_dataIn_E[58]
  PIN dyn2_dataIn_E[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END dyn2_dataIn_E[59]
  PIN dyn2_dataIn_E[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.330 0.000 2389.610 4.000 ;
    END
  END dyn2_dataIn_E[5]
  PIN dyn2_dataIn_E[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2315.440 2500.000 2316.040 ;
    END
  END dyn2_dataIn_E[60]
  PIN dyn2_dataIn_E[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.370 2496.000 2170.650 2500.000 ;
    END
  END dyn2_dataIn_E[61]
  PIN dyn2_dataIn_E[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END dyn2_dataIn_E[62]
  PIN dyn2_dataIn_E[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 2496.000 467.270 2500.000 ;
    END
  END dyn2_dataIn_E[63]
  PIN dyn2_dataIn_E[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 2496.000 1343.110 2500.000 ;
    END
  END dyn2_dataIn_E[6]
  PIN dyn2_dataIn_E[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 819.440 2500.000 820.040 ;
    END
  END dyn2_dataIn_E[7]
  PIN dyn2_dataIn_E[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2485.440 2500.000 2486.040 ;
    END
  END dyn2_dataIn_E[8]
  PIN dyn2_dataIn_E[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.170 2496.000 2299.450 2500.000 ;
    END
  END dyn2_dataIn_E[9]
  PIN dyn2_dataIn_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END dyn2_dataIn_N[0]
  PIN dyn2_dataIn_N[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 632.440 2500.000 633.040 ;
    END
  END dyn2_dataIn_N[10]
  PIN dyn2_dataIn_N[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.870 2496.000 2412.150 2500.000 ;
    END
  END dyn2_dataIn_N[11]
  PIN dyn2_dataIn_N[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2223.640 2500.000 2224.240 ;
    END
  END dyn2_dataIn_N[12]
  PIN dyn2_dataIn_N[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 2496.000 850.450 2500.000 ;
    END
  END dyn2_dataIn_N[13]
  PIN dyn2_dataIn_N[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 639.240 2500.000 639.840 ;
    END
  END dyn2_dataIn_N[14]
  PIN dyn2_dataIn_N[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 4.000 1850.240 ;
    END
  END dyn2_dataIn_N[15]
  PIN dyn2_dataIn_N[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1989.040 4.000 1989.640 ;
    END
  END dyn2_dataIn_N[16]
  PIN dyn2_dataIn_N[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END dyn2_dataIn_N[17]
  PIN dyn2_dataIn_N[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 2496.000 1001.790 2500.000 ;
    END
  END dyn2_dataIn_N[18]
  PIN dyn2_dataIn_N[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 4.000 ;
    END
  END dyn2_dataIn_N[19]
  PIN dyn2_dataIn_N[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1832.640 4.000 1833.240 ;
    END
  END dyn2_dataIn_N[1]
  PIN dyn2_dataIn_N[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 2496.000 1162.790 2500.000 ;
    END
  END dyn2_dataIn_N[20]
  PIN dyn2_dataIn_N[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1275.040 2500.000 1275.640 ;
    END
  END dyn2_dataIn_N[21]
  PIN dyn2_dataIn_N[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2155.640 2500.000 2156.240 ;
    END
  END dyn2_dataIn_N[22]
  PIN dyn2_dataIn_N[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1618.440 2500.000 1619.040 ;
    END
  END dyn2_dataIn_N[23]
  PIN dyn2_dataIn_N[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 2496.000 1191.770 2500.000 ;
    END
  END dyn2_dataIn_N[24]
  PIN dyn2_dataIn_N[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END dyn2_dataIn_N[25]
  PIN dyn2_dataIn_N[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 0.000 1246.510 4.000 ;
    END
  END dyn2_dataIn_N[26]
  PIN dyn2_dataIn_N[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1213.840 2500.000 1214.440 ;
    END
  END dyn2_dataIn_N[27]
  PIN dyn2_dataIn_N[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 0.000 1655.450 4.000 ;
    END
  END dyn2_dataIn_N[28]
  PIN dyn2_dataIn_N[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END dyn2_dataIn_N[29]
  PIN dyn2_dataIn_N[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END dyn2_dataIn_N[2]
  PIN dyn2_dataIn_N[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 2496.000 786.050 2500.000 ;
    END
  END dyn2_dataIn_N[30]
  PIN dyn2_dataIn_N[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END dyn2_dataIn_N[31]
  PIN dyn2_dataIn_N[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 231.240 2500.000 231.840 ;
    END
  END dyn2_dataIn_N[32]
  PIN dyn2_dataIn_N[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 2496.000 847.230 2500.000 ;
    END
  END dyn2_dataIn_N[33]
  PIN dyn2_dataIn_N[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 0.000 1494.450 4.000 ;
    END
  END dyn2_dataIn_N[34]
  PIN dyn2_dataIn_N[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.290 0.000 2286.570 4.000 ;
    END
  END dyn2_dataIn_N[35]
  PIN dyn2_dataIn_N[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 2496.000 1233.630 2500.000 ;
    END
  END dyn2_dataIn_N[36]
  PIN dyn2_dataIn_N[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2203.240 2500.000 2203.840 ;
    END
  END dyn2_dataIn_N[37]
  PIN dyn2_dataIn_N[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END dyn2_dataIn_N[38]
  PIN dyn2_dataIn_N[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2009.440 2500.000 2010.040 ;
    END
  END dyn2_dataIn_N[39]
  PIN dyn2_dataIn_N[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END dyn2_dataIn_N[3]
  PIN dyn2_dataIn_N[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1111.840 2500.000 1112.440 ;
    END
  END dyn2_dataIn_N[40]
  PIN dyn2_dataIn_N[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END dyn2_dataIn_N[41]
  PIN dyn2_dataIn_N[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2206.640 4.000 2207.240 ;
    END
  END dyn2_dataIn_N[42]
  PIN dyn2_dataIn_N[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 2496.000 1304.470 2500.000 ;
    END
  END dyn2_dataIn_N[43]
  PIN dyn2_dataIn_N[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2179.440 2500.000 2180.040 ;
    END
  END dyn2_dataIn_N[44]
  PIN dyn2_dataIn_N[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 2496.000 1281.930 2500.000 ;
    END
  END dyn2_dataIn_N[45]
  PIN dyn2_dataIn_N[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 2496.000 760.290 2500.000 ;
    END
  END dyn2_dataIn_N[46]
  PIN dyn2_dataIn_N[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2415.090 2496.000 2415.370 2500.000 ;
    END
  END dyn2_dataIn_N[47]
  PIN dyn2_dataIn_N[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END dyn2_dataIn_N[48]
  PIN dyn2_dataIn_N[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 2496.000 373.890 2500.000 ;
    END
  END dyn2_dataIn_N[49]
  PIN dyn2_dataIn_N[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END dyn2_dataIn_N[4]
  PIN dyn2_dataIn_N[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END dyn2_dataIn_N[50]
  PIN dyn2_dataIn_N[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END dyn2_dataIn_N[51]
  PIN dyn2_dataIn_N[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 2496.000 357.790 2500.000 ;
    END
  END dyn2_dataIn_N[52]
  PIN dyn2_dataIn_N[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END dyn2_dataIn_N[53]
  PIN dyn2_dataIn_N[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 40.840 2500.000 41.440 ;
    END
  END dyn2_dataIn_N[54]
  PIN dyn2_dataIn_N[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END dyn2_dataIn_N[55]
  PIN dyn2_dataIn_N[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 2496.000 753.850 2500.000 ;
    END
  END dyn2_dataIn_N[56]
  PIN dyn2_dataIn_N[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END dyn2_dataIn_N[57]
  PIN dyn2_dataIn_N[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 2496.000 1117.710 2500.000 ;
    END
  END dyn2_dataIn_N[58]
  PIN dyn2_dataIn_N[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1050.640 2500.000 1051.240 ;
    END
  END dyn2_dataIn_N[59]
  PIN dyn2_dataIn_N[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.130 2496.000 2196.410 2500.000 ;
    END
  END dyn2_dataIn_N[5]
  PIN dyn2_dataIn_N[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 2496.000 2270.470 2500.000 ;
    END
  END dyn2_dataIn_N[60]
  PIN dyn2_dataIn_N[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2471.840 4.000 2472.440 ;
    END
  END dyn2_dataIn_N[61]
  PIN dyn2_dataIn_N[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END dyn2_dataIn_N[62]
  PIN dyn2_dataIn_N[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.250 0.000 2344.530 4.000 ;
    END
  END dyn2_dataIn_N[63]
  PIN dyn2_dataIn_N[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 2496.000 505.910 2500.000 ;
    END
  END dyn2_dataIn_N[6]
  PIN dyn2_dataIn_N[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1227.440 2500.000 1228.040 ;
    END
  END dyn2_dataIn_N[7]
  PIN dyn2_dataIn_N[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END dyn2_dataIn_N[8]
  PIN dyn2_dataIn_N[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END dyn2_dataIn_N[9]
  PIN dyn2_dataIn_S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END dyn2_dataIn_S[0]
  PIN dyn2_dataIn_S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END dyn2_dataIn_S[10]
  PIN dyn2_dataIn_S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 493.040 2500.000 493.640 ;
    END
  END dyn2_dataIn_S[11]
  PIN dyn2_dataIn_S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.130 2496.000 2357.410 2500.000 ;
    END
  END dyn2_dataIn_S[12]
  PIN dyn2_dataIn_S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2441.240 2500.000 2441.840 ;
    END
  END dyn2_dataIn_S[13]
  PIN dyn2_dataIn_S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 2496.000 708.770 2500.000 ;
    END
  END dyn2_dataIn_S[14]
  PIN dyn2_dataIn_S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2414.040 4.000 2414.640 ;
    END
  END dyn2_dataIn_S[15]
  PIN dyn2_dataIn_S[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END dyn2_dataIn_S[16]
  PIN dyn2_dataIn_S[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END dyn2_dataIn_S[17]
  PIN dyn2_dataIn_S[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1669.440 4.000 1670.040 ;
    END
  END dyn2_dataIn_S[18]
  PIN dyn2_dataIn_S[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 972.440 2500.000 973.040 ;
    END
  END dyn2_dataIn_S[19]
  PIN dyn2_dataIn_S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END dyn2_dataIn_S[1]
  PIN dyn2_dataIn_S[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.210 2496.000 1919.490 2500.000 ;
    END
  END dyn2_dataIn_S[20]
  PIN dyn2_dataIn_S[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 2496.000 1565.290 2500.000 ;
    END
  END dyn2_dataIn_S[21]
  PIN dyn2_dataIn_S[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2274.640 4.000 2275.240 ;
    END
  END dyn2_dataIn_S[22]
  PIN dyn2_dataIn_S[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 105.440 2500.000 106.040 ;
    END
  END dyn2_dataIn_S[23]
  PIN dyn2_dataIn_S[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 2496.000 1642.570 2500.000 ;
    END
  END dyn2_dataIn_S[24]
  PIN dyn2_dataIn_S[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1394.040 2500.000 1394.640 ;
    END
  END dyn2_dataIn_S[25]
  PIN dyn2_dataIn_S[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END dyn2_dataIn_S[26]
  PIN dyn2_dataIn_S[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2142.040 2500.000 2142.640 ;
    END
  END dyn2_dataIn_S[27]
  PIN dyn2_dataIn_S[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END dyn2_dataIn_S[28]
  PIN dyn2_dataIn_S[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END dyn2_dataIn_S[29]
  PIN dyn2_dataIn_S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 2496.000 122.730 2500.000 ;
    END
  END dyn2_dataIn_S[2]
  PIN dyn2_dataIn_S[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 2496.000 2225.390 2500.000 ;
    END
  END dyn2_dataIn_S[30]
  PIN dyn2_dataIn_S[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END dyn2_dataIn_S[31]
  PIN dyn2_dataIn_S[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 2496.000 1665.110 2500.000 ;
    END
  END dyn2_dataIn_S[32]
  PIN dyn2_dataIn_S[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END dyn2_dataIn_S[33]
  PIN dyn2_dataIn_S[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END dyn2_dataIn_S[34]
  PIN dyn2_dataIn_S[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END dyn2_dataIn_S[35]
  PIN dyn2_dataIn_S[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END dyn2_dataIn_S[36]
  PIN dyn2_dataIn_S[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1353.240 2500.000 1353.840 ;
    END
  END dyn2_dataIn_S[37]
  PIN dyn2_dataIn_S[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 2496.000 2257.590 2500.000 ;
    END
  END dyn2_dataIn_S[38]
  PIN dyn2_dataIn_S[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 85.040 2500.000 85.640 ;
    END
  END dyn2_dataIn_S[39]
  PIN dyn2_dataIn_S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.970 0.000 1945.250 4.000 ;
    END
  END dyn2_dataIn_S[3]
  PIN dyn2_dataIn_S[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 2496.000 328.810 2500.000 ;
    END
  END dyn2_dataIn_S[40]
  PIN dyn2_dataIn_S[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 2496.000 538.110 2500.000 ;
    END
  END dyn2_dataIn_S[41]
  PIN dyn2_dataIn_S[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END dyn2_dataIn_S[42]
  PIN dyn2_dataIn_S[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2002.640 2500.000 2003.240 ;
    END
  END dyn2_dataIn_S[43]
  PIN dyn2_dataIn_S[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 374.040 2500.000 374.640 ;
    END
  END dyn2_dataIn_S[44]
  PIN dyn2_dataIn_S[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1499.440 4.000 1500.040 ;
    END
  END dyn2_dataIn_S[45]
  PIN dyn2_dataIn_S[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END dyn2_dataIn_S[46]
  PIN dyn2_dataIn_S[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 2496.000 1214.310 2500.000 ;
    END
  END dyn2_dataIn_S[47]
  PIN dyn2_dataIn_S[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1713.640 4.000 1714.240 ;
    END
  END dyn2_dataIn_S[48]
  PIN dyn2_dataIn_S[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END dyn2_dataIn_S[49]
  PIN dyn2_dataIn_S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.930 0.000 1681.210 4.000 ;
    END
  END dyn2_dataIn_S[4]
  PIN dyn2_dataIn_S[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END dyn2_dataIn_S[50]
  PIN dyn2_dataIn_S[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END dyn2_dataIn_S[51]
  PIN dyn2_dataIn_S[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.990 0.000 2238.270 4.000 ;
    END
  END dyn2_dataIn_S[52]
  PIN dyn2_dataIn_S[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 2496.000 959.930 2500.000 ;
    END
  END dyn2_dataIn_S[53]
  PIN dyn2_dataIn_S[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 462.440 2500.000 463.040 ;
    END
  END dyn2_dataIn_S[54]
  PIN dyn2_dataIn_S[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1696.640 2500.000 1697.240 ;
    END
  END dyn2_dataIn_S[55]
  PIN dyn2_dataIn_S[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END dyn2_dataIn_S[56]
  PIN dyn2_dataIn_S[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1934.640 4.000 1935.240 ;
    END
  END dyn2_dataIn_S[57]
  PIN dyn2_dataIn_S[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END dyn2_dataIn_S[58]
  PIN dyn2_dataIn_S[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.730 0.000 2132.010 4.000 ;
    END
  END dyn2_dataIn_S[59]
  PIN dyn2_dataIn_S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 2496.000 351.350 2500.000 ;
    END
  END dyn2_dataIn_S[5]
  PIN dyn2_dataIn_S[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END dyn2_dataIn_S[60]
  PIN dyn2_dataIn_S[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 421.640 2500.000 422.240 ;
    END
  END dyn2_dataIn_S[61]
  PIN dyn2_dataIn_S[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 13.640 2500.000 14.240 ;
    END
  END dyn2_dataIn_S[62]
  PIN dyn2_dataIn_S[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 2496.000 1690.870 2500.000 ;
    END
  END dyn2_dataIn_S[63]
  PIN dyn2_dataIn_S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END dyn2_dataIn_S[6]
  PIN dyn2_dataIn_S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 2496.000 1301.250 2500.000 ;
    END
  END dyn2_dataIn_S[7]
  PIN dyn2_dataIn_S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 2496.000 1243.290 2500.000 ;
    END
  END dyn2_dataIn_S[8]
  PIN dyn2_dataIn_S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 0.000 1797.130 4.000 ;
    END
  END dyn2_dataIn_S[9]
  PIN dyn2_dataIn_W[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 2496.000 1513.770 2500.000 ;
    END
  END dyn2_dataIn_W[0]
  PIN dyn2_dataIn_W[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2114.840 4.000 2115.440 ;
    END
  END dyn2_dataIn_W[10]
  PIN dyn2_dataIn_W[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2342.640 2500.000 2343.240 ;
    END
  END dyn2_dataIn_W[11]
  PIN dyn2_dataIn_W[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 2496.000 1597.490 2500.000 ;
    END
  END dyn2_dataIn_W[12]
  PIN dyn2_dataIn_W[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2230.440 4.000 2231.040 ;
    END
  END dyn2_dataIn_W[13]
  PIN dyn2_dataIn_W[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 2496.000 554.210 2500.000 ;
    END
  END dyn2_dataIn_W[14]
  PIN dyn2_dataIn_W[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END dyn2_dataIn_W[15]
  PIN dyn2_dataIn_W[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1611.640 2500.000 1612.240 ;
    END
  END dyn2_dataIn_W[16]
  PIN dyn2_dataIn_W[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 2496.000 972.810 2500.000 ;
    END
  END dyn2_dataIn_W[17]
  PIN dyn2_dataIn_W[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 438.640 2500.000 439.240 ;
    END
  END dyn2_dataIn_W[18]
  PIN dyn2_dataIn_W[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 0.000 1890.510 4.000 ;
    END
  END dyn2_dataIn_W[19]
  PIN dyn2_dataIn_W[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 2496.000 257.970 2500.000 ;
    END
  END dyn2_dataIn_W[1]
  PIN dyn2_dataIn_W[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END dyn2_dataIn_W[20]
  PIN dyn2_dataIn_W[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END dyn2_dataIn_W[21]
  PIN dyn2_dataIn_W[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END dyn2_dataIn_W[22]
  PIN dyn2_dataIn_W[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 918.040 2500.000 918.640 ;
    END
  END dyn2_dataIn_W[23]
  PIN dyn2_dataIn_W[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END dyn2_dataIn_W[24]
  PIN dyn2_dataIn_W[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 2496.000 1111.270 2500.000 ;
    END
  END dyn2_dataIn_W[25]
  PIN dyn2_dataIn_W[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2101.240 2500.000 2101.840 ;
    END
  END dyn2_dataIn_W[26]
  PIN dyn2_dataIn_W[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1135.640 2500.000 1136.240 ;
    END
  END dyn2_dataIn_W[27]
  PIN dyn2_dataIn_W[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END dyn2_dataIn_W[28]
  PIN dyn2_dataIn_W[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END dyn2_dataIn_W[29]
  PIN dyn2_dataIn_W[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END dyn2_dataIn_W[2]
  PIN dyn2_dataIn_W[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 2496.000 940.610 2500.000 ;
    END
  END dyn2_dataIn_W[30]
  PIN dyn2_dataIn_W[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END dyn2_dataIn_W[31]
  PIN dyn2_dataIn_W[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 969.040 2500.000 969.640 ;
    END
  END dyn2_dataIn_W[32]
  PIN dyn2_dataIn_W[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 2496.000 876.210 2500.000 ;
    END
  END dyn2_dataIn_W[33]
  PIN dyn2_dataIn_W[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.550 2496.000 1587.830 2500.000 ;
    END
  END dyn2_dataIn_W[34]
  PIN dyn2_dataIn_W[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END dyn2_dataIn_W[35]
  PIN dyn2_dataIn_W[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END dyn2_dataIn_W[36]
  PIN dyn2_dataIn_W[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1173.040 2500.000 1173.640 ;
    END
  END dyn2_dataIn_W[37]
  PIN dyn2_dataIn_W[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 2496.000 1062.970 2500.000 ;
    END
  END dyn2_dataIn_W[38]
  PIN dyn2_dataIn_W[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 2496.000 534.890 2500.000 ;
    END
  END dyn2_dataIn_W[39]
  PIN dyn2_dataIn_W[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END dyn2_dataIn_W[3]
  PIN dyn2_dataIn_W[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2448.040 4.000 2448.640 ;
    END
  END dyn2_dataIn_W[40]
  PIN dyn2_dataIn_W[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 2496.000 435.070 2500.000 ;
    END
  END dyn2_dataIn_W[41]
  PIN dyn2_dataIn_W[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 360.440 2500.000 361.040 ;
    END
  END dyn2_dataIn_W[42]
  PIN dyn2_dataIn_W[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.040 4.000 935.640 ;
    END
  END dyn2_dataIn_W[43]
  PIN dyn2_dataIn_W[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END dyn2_dataIn_W[44]
  PIN dyn2_dataIn_W[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.030 2496.000 1697.310 2500.000 ;
    END
  END dyn2_dataIn_W[45]
  PIN dyn2_dataIn_W[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END dyn2_dataIn_W[46]
  PIN dyn2_dataIn_W[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 0.000 1864.750 4.000 ;
    END
  END dyn2_dataIn_W[47]
  PIN dyn2_dataIn_W[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END dyn2_dataIn_W[48]
  PIN dyn2_dataIn_W[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.510 0.000 2450.790 4.000 ;
    END
  END dyn2_dataIn_W[49]
  PIN dyn2_dataIn_W[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 2496.000 325.590 2500.000 ;
    END
  END dyn2_dataIn_W[4]
  PIN dyn2_dataIn_W[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 2496.000 386.770 2500.000 ;
    END
  END dyn2_dataIn_W[50]
  PIN dyn2_dataIn_W[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END dyn2_dataIn_W[51]
  PIN dyn2_dataIn_W[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1397.440 2500.000 1398.040 ;
    END
  END dyn2_dataIn_W[52]
  PIN dyn2_dataIn_W[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2077.440 2500.000 2078.040 ;
    END
  END dyn2_dataIn_W[53]
  PIN dyn2_dataIn_W[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END dyn2_dataIn_W[54]
  PIN dyn2_dataIn_W[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.710 2496.000 2482.990 2500.000 ;
    END
  END dyn2_dataIn_W[55]
  PIN dyn2_dataIn_W[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1863.240 2500.000 1863.840 ;
    END
  END dyn2_dataIn_W[56]
  PIN dyn2_dataIn_W[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END dyn2_dataIn_W[57]
  PIN dyn2_dataIn_W[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1880.240 4.000 1880.840 ;
    END
  END dyn2_dataIn_W[58]
  PIN dyn2_dataIn_W[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END dyn2_dataIn_W[59]
  PIN dyn2_dataIn_W[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END dyn2_dataIn_W[5]
  PIN dyn2_dataIn_W[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2199.840 4.000 2200.440 ;
    END
  END dyn2_dataIn_W[60]
  PIN dyn2_dataIn_W[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 2496.000 148.490 2500.000 ;
    END
  END dyn2_dataIn_W[61]
  PIN dyn2_dataIn_W[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1336.240 2500.000 1336.840 ;
    END
  END dyn2_dataIn_W[62]
  PIN dyn2_dataIn_W[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 622.240 2500.000 622.840 ;
    END
  END dyn2_dataIn_W[63]
  PIN dyn2_dataIn_W[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 183.640 2500.000 184.240 ;
    END
  END dyn2_dataIn_W[6]
  PIN dyn2_dataIn_W[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END dyn2_dataIn_W[7]
  PIN dyn2_dataIn_W[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END dyn2_dataIn_W[8]
  PIN dyn2_dataIn_W[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 795.640 2500.000 796.240 ;
    END
  END dyn2_dataIn_W[9]
  PIN dyn2_validIn_E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 394.440 2500.000 395.040 ;
    END
  END dyn2_validIn_E
  PIN dyn2_validIn_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END dyn2_validIn_N
  PIN dyn2_validIn_S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END dyn2_validIn_S
  PIN dyn2_validIn_W
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 2496.000 637.930 2500.000 ;
    END
  END dyn2_validIn_W
  PIN dyn2_yummyOut_E
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END dyn2_yummyOut_E
  PIN dyn2_yummyOut_N
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 326.440 2500.000 327.040 ;
    END
  END dyn2_yummyOut_N
  PIN dyn2_yummyOut_S
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 2496.000 460.830 2500.000 ;
    END
  END dyn2_yummyOut_S
  PIN dyn2_yummyOut_W
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END dyn2_yummyOut_W
  PIN flat_tileid[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END flat_tileid[0]
  PIN flat_tileid[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.790 2496.000 2206.070 2500.000 ;
    END
  END flat_tileid[1]
  PIN flat_tileid[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2492.240 4.000 2492.840 ;
    END
  END flat_tileid[2]
  PIN flat_tileid[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2016.240 4.000 2016.840 ;
    END
  END flat_tileid[3]
  PIN flat_tileid[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2335.840 2500.000 2336.440 ;
    END
  END flat_tileid[4]
  PIN flat_tileid[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 0.040 2500.000 0.640 ;
    END
  END flat_tileid[5]
  PIN flat_tileid[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.370 0.000 2331.650 4.000 ;
    END
  END flat_tileid[6]
  PIN flat_tileid[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.250 2496.000 2344.530 2500.000 ;
    END
  END flat_tileid[7]
  PIN jtag_tiles_ucb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 2496.000 48.670 2500.000 ;
    END
  END jtag_tiles_ucb_data[0]
  PIN jtag_tiles_ucb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 2496.000 789.270 2500.000 ;
    END
  END jtag_tiles_ucb_data[1]
  PIN jtag_tiles_ucb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2087.640 4.000 2088.240 ;
    END
  END jtag_tiles_ucb_data[2]
  PIN jtag_tiles_ucb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 2496.000 1040.430 2500.000 ;
    END
  END jtag_tiles_ucb_data[3]
  PIN jtag_tiles_ucb_val
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 0.000 1578.170 4.000 ;
    END
  END jtag_tiles_ucb_val
  PIN l15_config_req_address_s2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 2496.000 1932.370 2500.000 ;
    END
  END l15_config_req_address_s2[10]
  PIN l15_config_req_address_s2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 2496.000 1481.570 2500.000 ;
    END
  END l15_config_req_address_s2[11]
  PIN l15_config_req_address_s2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END l15_config_req_address_s2[12]
  PIN l15_config_req_address_s2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.770 2496.000 1591.050 2500.000 ;
    END
  END l15_config_req_address_s2[13]
  PIN l15_config_req_address_s2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 3.440 2500.000 4.040 ;
    END
  END l15_config_req_address_s2[14]
  PIN l15_config_req_address_s2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1475.640 2500.000 1476.240 ;
    END
  END l15_config_req_address_s2[15]
  PIN l15_config_req_address_s2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2305.240 4.000 2305.840 ;
    END
  END l15_config_req_address_s2[8]
  PIN l15_config_req_address_s2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END l15_config_req_address_s2[9]
  PIN l15_config_req_rw_s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 2496.000 615.390 2500.000 ;
    END
  END l15_config_req_rw_s2
  PIN l15_config_req_val_s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 999.640 2500.000 1000.240 ;
    END
  END l15_config_req_val_s2
  PIN l15_config_write_req_data_s2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END l15_config_write_req_data_s2[0]
  PIN l15_config_write_req_data_s2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END l15_config_write_req_data_s2[10]
  PIN l15_config_write_req_data_s2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2376.640 2500.000 2377.240 ;
    END
  END l15_config_write_req_data_s2[11]
  PIN l15_config_write_req_data_s2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 2496.000 1362.430 2500.000 ;
    END
  END l15_config_write_req_data_s2[12]
  PIN l15_config_write_req_data_s2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 2496.000 1835.770 2500.000 ;
    END
  END l15_config_write_req_data_s2[13]
  PIN l15_config_write_req_data_s2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 180.240 2500.000 180.840 ;
    END
  END l15_config_write_req_data_s2[14]
  PIN l15_config_write_req_data_s2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END l15_config_write_req_data_s2[15]
  PIN l15_config_write_req_data_s2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 0.000 1500.890 4.000 ;
    END
  END l15_config_write_req_data_s2[16]
  PIN l15_config_write_req_data_s2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2356.240 2500.000 2356.840 ;
    END
  END l15_config_write_req_data_s2[17]
  PIN l15_config_write_req_data_s2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 397.840 2500.000 398.440 ;
    END
  END l15_config_write_req_data_s2[18]
  PIN l15_config_write_req_data_s2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END l15_config_write_req_data_s2[19]
  PIN l15_config_write_req_data_s2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 2496.000 1703.750 2500.000 ;
    END
  END l15_config_write_req_data_s2[1]
  PIN l15_config_write_req_data_s2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2420.840 4.000 2421.440 ;
    END
  END l15_config_write_req_data_s2[20]
  PIN l15_config_write_req_data_s2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1924.440 4.000 1925.040 ;
    END
  END l15_config_write_req_data_s2[21]
  PIN l15_config_write_req_data_s2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1778.240 2500.000 1778.840 ;
    END
  END l15_config_write_req_data_s2[22]
  PIN l15_config_write_req_data_s2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END l15_config_write_req_data_s2[23]
  PIN l15_config_write_req_data_s2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 2496.000 512.350 2500.000 ;
    END
  END l15_config_write_req_data_s2[24]
  PIN l15_config_write_req_data_s2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2281.440 2500.000 2282.040 ;
    END
  END l15_config_write_req_data_s2[25]
  PIN l15_config_write_req_data_s2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END l15_config_write_req_data_s2[26]
  PIN l15_config_write_req_data_s2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 2496.000 792.490 2500.000 ;
    END
  END l15_config_write_req_data_s2[27]
  PIN l15_config_write_req_data_s2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END l15_config_write_req_data_s2[28]
  PIN l15_config_write_req_data_s2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2495.640 4.000 2496.240 ;
    END
  END l15_config_write_req_data_s2[29]
  PIN l15_config_write_req_data_s2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.890 0.000 2383.170 4.000 ;
    END
  END l15_config_write_req_data_s2[2]
  PIN l15_config_write_req_data_s2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1278.440 2500.000 1279.040 ;
    END
  END l15_config_write_req_data_s2[30]
  PIN l15_config_write_req_data_s2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 2496.000 1330.230 2500.000 ;
    END
  END l15_config_write_req_data_s2[31]
  PIN l15_config_write_req_data_s2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 2496.000 2354.190 2500.000 ;
    END
  END l15_config_write_req_data_s2[32]
  PIN l15_config_write_req_data_s2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END l15_config_write_req_data_s2[33]
  PIN l15_config_write_req_data_s2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END l15_config_write_req_data_s2[34]
  PIN l15_config_write_req_data_s2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1315.840 2500.000 1316.440 ;
    END
  END l15_config_write_req_data_s2[35]
  PIN l15_config_write_req_data_s2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 2496.000 576.750 2500.000 ;
    END
  END l15_config_write_req_data_s2[36]
  PIN l15_config_write_req_data_s2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END l15_config_write_req_data_s2[37]
  PIN l15_config_write_req_data_s2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 2496.000 431.850 2500.000 ;
    END
  END l15_config_write_req_data_s2[38]
  PIN l15_config_write_req_data_s2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 921.440 2500.000 922.040 ;
    END
  END l15_config_write_req_data_s2[39]
  PIN l15_config_write_req_data_s2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 2496.000 1005.010 2500.000 ;
    END
  END l15_config_write_req_data_s2[3]
  PIN l15_config_write_req_data_s2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END l15_config_write_req_data_s2[40]
  PIN l15_config_write_req_data_s2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END l15_config_write_req_data_s2[41]
  PIN l15_config_write_req_data_s2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END l15_config_write_req_data_s2[42]
  PIN l15_config_write_req_data_s2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END l15_config_write_req_data_s2[43]
  PIN l15_config_write_req_data_s2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 2496.000 1948.470 2500.000 ;
    END
  END l15_config_write_req_data_s2[44]
  PIN l15_config_write_req_data_s2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 2496.000 882.650 2500.000 ;
    END
  END l15_config_write_req_data_s2[45]
  PIN l15_config_write_req_data_s2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 2496.000 315.930 2500.000 ;
    END
  END l15_config_write_req_data_s2[46]
  PIN l15_config_write_req_data_s2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 0.000 1459.030 4.000 ;
    END
  END l15_config_write_req_data_s2[47]
  PIN l15_config_write_req_data_s2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2237.240 2500.000 2237.840 ;
    END
  END l15_config_write_req_data_s2[48]
  PIN l15_config_write_req_data_s2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1373.640 2500.000 1374.240 ;
    END
  END l15_config_write_req_data_s2[49]
  PIN l15_config_write_req_data_s2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END l15_config_write_req_data_s2[4]
  PIN l15_config_write_req_data_s2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2322.240 4.000 2322.840 ;
    END
  END l15_config_write_req_data_s2[50]
  PIN l15_config_write_req_data_s2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1805.440 4.000 1806.040 ;
    END
  END l15_config_write_req_data_s2[51]
  PIN l15_config_write_req_data_s2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END l15_config_write_req_data_s2[52]
  PIN l15_config_write_req_data_s2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 618.840 2500.000 619.440 ;
    END
  END l15_config_write_req_data_s2[53]
  PIN l15_config_write_req_data_s2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END l15_config_write_req_data_s2[54]
  PIN l15_config_write_req_data_s2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END l15_config_write_req_data_s2[55]
  PIN l15_config_write_req_data_s2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 948.640 2500.000 949.240 ;
    END
  END l15_config_write_req_data_s2[56]
  PIN l15_config_write_req_data_s2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1536.840 2500.000 1537.440 ;
    END
  END l15_config_write_req_data_s2[57]
  PIN l15_config_write_req_data_s2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 873.840 2500.000 874.440 ;
    END
  END l15_config_write_req_data_s2[58]
  PIN l15_config_write_req_data_s2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 2496.000 802.150 2500.000 ;
    END
  END l15_config_write_req_data_s2[59]
  PIN l15_config_write_req_data_s2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2298.440 2500.000 2299.040 ;
    END
  END l15_config_write_req_data_s2[5]
  PIN l15_config_write_req_data_s2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END l15_config_write_req_data_s2[60]
  PIN l15_config_write_req_data_s2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 2496.000 750.630 2500.000 ;
    END
  END l15_config_write_req_data_s2[61]
  PIN l15_config_write_req_data_s2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END l15_config_write_req_data_s2[62]
  PIN l15_config_write_req_data_s2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.730 0.000 2454.010 4.000 ;
    END
  END l15_config_write_req_data_s2[63]
  PIN l15_config_write_req_data_s2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END l15_config_write_req_data_s2[6]
  PIN l15_config_write_req_data_s2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END l15_config_write_req_data_s2[7]
  PIN l15_config_write_req_data_s2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END l15_config_write_req_data_s2[8]
  PIN l15_config_write_req_data_s2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 2496.000 718.430 2500.000 ;
    END
  END l15_config_write_req_data_s2[9]
  PIN l15_dmbr_l1missIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END l15_dmbr_l1missIn
  PIN l15_dmbr_l1missTag[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END l15_dmbr_l1missTag[0]
  PIN l15_dmbr_l1missTag[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 210.840 2500.000 211.440 ;
    END
  END l15_dmbr_l1missTag[1]
  PIN l15_dmbr_l1missTag[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END l15_dmbr_l1missTag[2]
  PIN l15_dmbr_l1missTag[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END l15_dmbr_l1missTag[3]
  PIN l15_dmbr_l2missIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 0.000 2070.830 4.000 ;
    END
  END l15_dmbr_l2missIn
  PIN l15_dmbr_l2missTag[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END l15_dmbr_l2missTag[0]
  PIN l15_dmbr_l2missTag[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 2496.000 177.470 2500.000 ;
    END
  END l15_dmbr_l2missTag[1]
  PIN l15_dmbr_l2missTag[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 2496.000 1610.370 2500.000 ;
    END
  END l15_dmbr_l2missTag[2]
  PIN l15_dmbr_l2missTag[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1013.240 2500.000 1013.840 ;
    END
  END l15_dmbr_l2missTag[3]
  PIN l15_dmbr_l2responseIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1077.840 2500.000 1078.440 ;
    END
  END l15_dmbr_l2responseIn
  PIN l15_transducer_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1295.440 2500.000 1296.040 ;
    END
  END l15_transducer_ack
  PIN l15_transducer_atomic
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 2496.000 1069.410 2500.000 ;
    END
  END l15_transducer_atomic
  PIN l15_transducer_blockinitstore
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END l15_transducer_blockinitstore
  PIN l15_transducer_cross_invalidate
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END l15_transducer_cross_invalidate
  PIN l15_transducer_cross_invalidate_way[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END l15_transducer_cross_invalidate_way[0]
  PIN l15_transducer_cross_invalidate_way[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.090 2496.000 2093.370 2500.000 ;
    END
  END l15_transducer_cross_invalidate_way[1]
  PIN l15_transducer_data_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.690 2496.000 2189.970 2500.000 ;
    END
  END l15_transducer_data_0[0]
  PIN l15_transducer_data_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 2496.000 2112.690 2500.000 ;
    END
  END l15_transducer_data_0[10]
  PIN l15_transducer_data_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2386.840 2500.000 2387.440 ;
    END
  END l15_transducer_data_0[11]
  PIN l15_transducer_data_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 533.840 2500.000 534.440 ;
    END
  END l15_transducer_data_0[12]
  PIN l15_transducer_data_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END l15_transducer_data_0[13]
  PIN l15_transducer_data_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 2496.000 1346.330 2500.000 ;
    END
  END l15_transducer_data_0[14]
  PIN l15_transducer_data_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1523.240 2500.000 1523.840 ;
    END
  END l15_transducer_data_0[15]
  PIN l15_transducer_data_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 2496.000 831.130 2500.000 ;
    END
  END l15_transducer_data_0[16]
  PIN l15_transducer_data_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1424.640 4.000 1425.240 ;
    END
  END l15_transducer_data_0[17]
  PIN l15_transducer_data_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.550 0.000 2392.830 4.000 ;
    END
  END l15_transducer_data_0[18]
  PIN l15_transducer_data_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END l15_transducer_data_0[19]
  PIN l15_transducer_data_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END l15_transducer_data_0[1]
  PIN l15_transducer_data_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END l15_transducer_data_0[20]
  PIN l15_transducer_data_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 125.840 2500.000 126.440 ;
    END
  END l15_transducer_data_0[21]
  PIN l15_transducer_data_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END l15_transducer_data_0[22]
  PIN l15_transducer_data_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 428.440 2500.000 429.040 ;
    END
  END l15_transducer_data_0[23]
  PIN l15_transducer_data_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.010 2496.000 2209.290 2500.000 ;
    END
  END l15_transducer_data_0[24]
  PIN l15_transducer_data_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END l15_transducer_data_0[25]
  PIN l15_transducer_data_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1652.440 2500.000 1653.040 ;
    END
  END l15_transducer_data_0[26]
  PIN l15_transducer_data_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 2496.000 1668.330 2500.000 ;
    END
  END l15_transducer_data_0[27]
  PIN l15_transducer_data_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1601.440 2500.000 1602.040 ;
    END
  END l15_transducer_data_0[28]
  PIN l15_transducer_data_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.890 2496.000 2061.170 2500.000 ;
    END
  END l15_transducer_data_0[29]
  PIN l15_transducer_data_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 520.240 2500.000 520.840 ;
    END
  END l15_transducer_data_0[2]
  PIN l15_transducer_data_0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END l15_transducer_data_0[30]
  PIN l15_transducer_data_0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2356.240 4.000 2356.840 ;
    END
  END l15_transducer_data_0[31]
  PIN l15_transducer_data_0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END l15_transducer_data_0[32]
  PIN l15_transducer_data_0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 2496.000 509.130 2500.000 ;
    END
  END l15_transducer_data_0[33]
  PIN l15_transducer_data_0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 2496.000 1671.550 2500.000 ;
    END
  END l15_transducer_data_0[34]
  PIN l15_transducer_data_0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 486.240 2500.000 486.840 ;
    END
  END l15_transducer_data_0[35]
  PIN l15_transducer_data_0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END l15_transducer_data_0[36]
  PIN l15_transducer_data_0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END l15_transducer_data_0[37]
  PIN l15_transducer_data_0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END l15_transducer_data_0[38]
  PIN l15_transducer_data_0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 2496.000 711.990 2500.000 ;
    END
  END l15_transducer_data_0[39]
  PIN l15_transducer_data_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2084.240 2500.000 2084.840 ;
    END
  END l15_transducer_data_0[3]
  PIN l15_transducer_data_0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.490 0.000 2479.770 4.000 ;
    END
  END l15_transducer_data_0[40]
  PIN l15_transducer_data_0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.650 2496.000 2408.930 2500.000 ;
    END
  END l15_transducer_data_0[41]
  PIN l15_transducer_data_0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.410 2496.000 2434.690 2500.000 ;
    END
  END l15_transducer_data_0[42]
  PIN l15_transducer_data_0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.040 4.000 1496.640 ;
    END
  END l15_transducer_data_0[43]
  PIN l15_transducer_data_0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1094.840 2500.000 1095.440 ;
    END
  END l15_transducer_data_0[44]
  PIN l15_transducer_data_0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.370 0.000 2009.650 4.000 ;
    END
  END l15_transducer_data_0[45]
  PIN l15_transducer_data_0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 0.000 1858.310 4.000 ;
    END
  END l15_transducer_data_0[46]
  PIN l15_transducer_data_0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END l15_transducer_data_0[47]
  PIN l15_transducer_data_0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 0.000 2431.470 4.000 ;
    END
  END l15_transducer_data_0[48]
  PIN l15_transducer_data_0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END l15_transducer_data_0[49]
  PIN l15_transducer_data_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2495.590 2496.000 2495.870 2500.000 ;
    END
  END l15_transducer_data_0[4]
  PIN l15_transducer_data_0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 2496.000 1327.010 2500.000 ;
    END
  END l15_transducer_data_0[50]
  PIN l15_transducer_data_0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END l15_transducer_data_0[51]
  PIN l15_transducer_data_0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.070 0.000 2283.350 4.000 ;
    END
  END l15_transducer_data_0[52]
  PIN l15_transducer_data_0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END l15_transducer_data_0[53]
  PIN l15_transducer_data_0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END l15_transducer_data_0[54]
  PIN l15_transducer_data_0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2415.090 0.000 2415.370 4.000 ;
    END
  END l15_transducer_data_0[55]
  PIN l15_transducer_data_0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2469.830 2496.000 2470.110 2500.000 ;
    END
  END l15_transducer_data_0[56]
  PIN l15_transducer_data_0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2043.440 2500.000 2044.040 ;
    END
  END l15_transducer_data_0[57]
  PIN l15_transducer_data_0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END l15_transducer_data_0[58]
  PIN l15_transducer_data_0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2070.640 4.000 2071.240 ;
    END
  END l15_transducer_data_0[59]
  PIN l15_transducer_data_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END l15_transducer_data_0[5]
  PIN l15_transducer_data_0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END l15_transducer_data_0[60]
  PIN l15_transducer_data_0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2220.240 4.000 2220.840 ;
    END
  END l15_transducer_data_0[61]
  PIN l15_transducer_data_0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 0.000 1542.750 4.000 ;
    END
  END l15_transducer_data_0[62]
  PIN l15_transducer_data_0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END l15_transducer_data_0[63]
  PIN l15_transducer_data_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.950 0.000 1974.230 4.000 ;
    END
  END l15_transducer_data_0[6]
  PIN l15_transducer_data_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END l15_transducer_data_0[7]
  PIN l15_transducer_data_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2182.840 4.000 2183.440 ;
    END
  END l15_transducer_data_0[8]
  PIN l15_transducer_data_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 2496.000 834.350 2500.000 ;
    END
  END l15_transducer_data_0[9]
  PIN l15_transducer_data_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2325.640 2500.000 2326.240 ;
    END
  END l15_transducer_data_1[0]
  PIN l15_transducer_data_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 2496.000 425.410 2500.000 ;
    END
  END l15_transducer_data_1[10]
  PIN l15_transducer_data_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 2496.000 1442.930 2500.000 ;
    END
  END l15_transducer_data_1[11]
  PIN l15_transducer_data_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END l15_transducer_data_1[12]
  PIN l15_transducer_data_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2138.640 2500.000 2139.240 ;
    END
  END l15_transducer_data_1[13]
  PIN l15_transducer_data_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END l15_transducer_data_1[14]
  PIN l15_transducer_data_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 2496.000 1430.050 2500.000 ;
    END
  END l15_transducer_data_1[15]
  PIN l15_transducer_data_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1533.440 2500.000 1534.040 ;
    END
  END l15_transducer_data_1[16]
  PIN l15_transducer_data_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END l15_transducer_data_1[17]
  PIN l15_transducer_data_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 863.640 2500.000 864.240 ;
    END
  END l15_transducer_data_1[18]
  PIN l15_transducer_data_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END l15_transducer_data_1[19]
  PIN l15_transducer_data_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2288.240 2500.000 2288.840 ;
    END
  END l15_transducer_data_1[1]
  PIN l15_transducer_data_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1754.440 2500.000 1755.040 ;
    END
  END l15_transducer_data_1[20]
  PIN l15_transducer_data_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 336.640 2500.000 337.240 ;
    END
  END l15_transducer_data_1[21]
  PIN l15_transducer_data_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.290 2496.000 2447.570 2500.000 ;
    END
  END l15_transducer_data_1[22]
  PIN l15_transducer_data_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1774.840 2500.000 1775.440 ;
    END
  END l15_transducer_data_1[23]
  PIN l15_transducer_data_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END l15_transducer_data_1[24]
  PIN l15_transducer_data_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 2496.000 525.230 2500.000 ;
    END
  END l15_transducer_data_1[25]
  PIN l15_transducer_data_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2250.840 2500.000 2251.440 ;
    END
  END l15_transducer_data_1[26]
  PIN l15_transducer_data_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1866.640 2500.000 1867.240 ;
    END
  END l15_transducer_data_1[27]
  PIN l15_transducer_data_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 2496.000 1046.870 2500.000 ;
    END
  END l15_transducer_data_1[28]
  PIN l15_transducer_data_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2264.440 4.000 2265.040 ;
    END
  END l15_transducer_data_1[29]
  PIN l15_transducer_data_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 2496.000 480.150 2500.000 ;
    END
  END l15_transducer_data_1[2]
  PIN l15_transducer_data_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2308.640 2500.000 2309.240 ;
    END
  END l15_transducer_data_1[30]
  PIN l15_transducer_data_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 2496.000 476.930 2500.000 ;
    END
  END l15_transducer_data_1[31]
  PIN l15_transducer_data_1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END l15_transducer_data_1[32]
  PIN l15_transducer_data_1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2063.840 4.000 2064.440 ;
    END
  END l15_transducer_data_1[33]
  PIN l15_transducer_data_1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 4.000 ;
    END
  END l15_transducer_data_1[34]
  PIN l15_transducer_data_1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2366.790 2496.000 2367.070 2500.000 ;
    END
  END l15_transducer_data_1[35]
  PIN l15_transducer_data_1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2451.440 2500.000 2452.040 ;
    END
  END l15_transducer_data_1[36]
  PIN l15_transducer_data_1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1530.040 2500.000 1530.640 ;
    END
  END l15_transducer_data_1[37]
  PIN l15_transducer_data_1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 2496.000 1095.170 2500.000 ;
    END
  END l15_transducer_data_1[38]
  PIN l15_transducer_data_1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1234.240 2500.000 1234.840 ;
    END
  END l15_transducer_data_1[39]
  PIN l15_transducer_data_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1251.240 2500.000 1251.840 ;
    END
  END l15_transducer_data_1[3]
  PIN l15_transducer_data_1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END l15_transducer_data_1[40]
  PIN l15_transducer_data_1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2210.040 2500.000 2210.640 ;
    END
  END l15_transducer_data_1[41]
  PIN l15_transducer_data_1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END l15_transducer_data_1[42]
  PIN l15_transducer_data_1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 261.840 2500.000 262.440 ;
    END
  END l15_transducer_data_1[43]
  PIN l15_transducer_data_1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 4.000 ;
    END
  END l15_transducer_data_1[44]
  PIN l15_transducer_data_1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END l15_transducer_data_1[45]
  PIN l15_transducer_data_1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END l15_transducer_data_1[46]
  PIN l15_transducer_data_1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2295.040 2500.000 2295.640 ;
    END
  END l15_transducer_data_1[47]
  PIN l15_transducer_data_1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 2496.000 380.330 2500.000 ;
    END
  END l15_transducer_data_1[48]
  PIN l15_transducer_data_1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2148.840 2500.000 2149.440 ;
    END
  END l15_transducer_data_1[49]
  PIN l15_transducer_data_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2386.840 4.000 2387.440 ;
    END
  END l15_transducer_data_1[4]
  PIN l15_transducer_data_1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END l15_transducer_data_1[50]
  PIN l15_transducer_data_1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2420.840 2500.000 2421.440 ;
    END
  END l15_transducer_data_1[51]
  PIN l15_transducer_data_1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 737.840 2500.000 738.440 ;
    END
  END l15_transducer_data_1[52]
  PIN l15_transducer_data_1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 979.240 2500.000 979.840 ;
    END
  END l15_transducer_data_1[53]
  PIN l15_transducer_data_1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 4.000 ;
    END
  END l15_transducer_data_1[54]
  PIN l15_transducer_data_1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 57.840 2500.000 58.440 ;
    END
  END l15_transducer_data_1[55]
  PIN l15_transducer_data_1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1054.040 2500.000 1054.640 ;
    END
  END l15_transducer_data_1[56]
  PIN l15_transducer_data_1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 2496.000 1401.070 2500.000 ;
    END
  END l15_transducer_data_1[57]
  PIN l15_transducer_data_1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1196.840 2500.000 1197.440 ;
    END
  END l15_transducer_data_1[58]
  PIN l15_transducer_data_1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END l15_transducer_data_1[59]
  PIN l15_transducer_data_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END l15_transducer_data_1[5]
  PIN l15_transducer_data_1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END l15_transducer_data_1[60]
  PIN l15_transducer_data_1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1071.040 2500.000 1071.640 ;
    END
  END l15_transducer_data_1[61]
  PIN l15_transducer_data_1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 4.000 ;
    END
  END l15_transducer_data_1[62]
  PIN l15_transducer_data_1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 2496.000 2148.110 2500.000 ;
    END
  END l15_transducer_data_1[63]
  PIN l15_transducer_data_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 2496.000 96.970 2500.000 ;
    END
  END l15_transducer_data_1[6]
  PIN l15_transducer_data_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 2496.000 1011.450 2500.000 ;
    END
  END l15_transducer_data_1[7]
  PIN l15_transducer_data_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1955.040 4.000 1955.640 ;
    END
  END l15_transducer_data_1[8]
  PIN l15_transducer_data_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END l15_transducer_data_1[9]
  PIN l15_transducer_data_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END l15_transducer_data_2[0]
  PIN l15_transducer_data_2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END l15_transducer_data_2[10]
  PIN l15_transducer_data_2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END l15_transducer_data_2[11]
  PIN l15_transducer_data_2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END l15_transducer_data_2[12]
  PIN l15_transducer_data_2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 47.640 2500.000 48.240 ;
    END
  END l15_transducer_data_2[13]
  PIN l15_transducer_data_2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END l15_transducer_data_2[14]
  PIN l15_transducer_data_2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END l15_transducer_data_2[15]
  PIN l15_transducer_data_2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 2496.000 1713.410 2500.000 ;
    END
  END l15_transducer_data_2[16]
  PIN l15_transducer_data_2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END l15_transducer_data_2[17]
  PIN l15_transducer_data_2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 163.240 2500.000 163.840 ;
    END
  END l15_transducer_data_2[18]
  PIN l15_transducer_data_2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1825.840 2500.000 1826.440 ;
    END
  END l15_transducer_data_2[19]
  PIN l15_transducer_data_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 0.000 1851.870 4.000 ;
    END
  END l15_transducer_data_2[1]
  PIN l15_transducer_data_2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END l15_transducer_data_2[20]
  PIN l15_transducer_data_2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 673.240 2500.000 673.840 ;
    END
  END l15_transducer_data_2[21]
  PIN l15_transducer_data_2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 2496.000 1903.390 2500.000 ;
    END
  END l15_transducer_data_2[22]
  PIN l15_transducer_data_2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2097.840 4.000 2098.440 ;
    END
  END l15_transducer_data_2[23]
  PIN l15_transducer_data_2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 805.840 2500.000 806.440 ;
    END
  END l15_transducer_data_2[24]
  PIN l15_transducer_data_2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1747.640 2500.000 1748.240 ;
    END
  END l15_transducer_data_2[25]
  PIN l15_transducer_data_2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.850 2496.000 2441.130 2500.000 ;
    END
  END l15_transducer_data_2[26]
  PIN l15_transducer_data_2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 2496.000 1829.330 2500.000 ;
    END
  END l15_transducer_data_2[27]
  PIN l15_transducer_data_2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1842.840 4.000 1843.440 ;
    END
  END l15_transducer_data_2[28]
  PIN l15_transducer_data_2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 2496.000 196.790 2500.000 ;
    END
  END l15_transducer_data_2[29]
  PIN l15_transducer_data_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END l15_transducer_data_2[2]
  PIN l15_transducer_data_2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END l15_transducer_data_2[30]
  PIN l15_transducer_data_2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1696.640 4.000 1697.240 ;
    END
  END l15_transducer_data_2[31]
  PIN l15_transducer_data_2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.210 2496.000 2402.490 2500.000 ;
    END
  END l15_transducer_data_2[32]
  PIN l15_transducer_data_2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END l15_transducer_data_2[33]
  PIN l15_transducer_data_2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END l15_transducer_data_2[34]
  PIN l15_transducer_data_2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END l15_transducer_data_2[35]
  PIN l15_transducer_data_2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2193.040 4.000 2193.640 ;
    END
  END l15_transducer_data_2[36]
  PIN l15_transducer_data_2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END l15_transducer_data_2[37]
  PIN l15_transducer_data_2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 0.000 1887.290 4.000 ;
    END
  END l15_transducer_data_2[38]
  PIN l15_transducer_data_2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1744.240 4.000 1744.840 ;
    END
  END l15_transducer_data_2[39]
  PIN l15_transducer_data_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END l15_transducer_data_2[3]
  PIN l15_transducer_data_2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 2496.000 454.390 2500.000 ;
    END
  END l15_transducer_data_2[40]
  PIN l15_transducer_data_2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END l15_transducer_data_2[41]
  PIN l15_transducer_data_2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END l15_transducer_data_2[42]
  PIN l15_transducer_data_2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 625.640 2500.000 626.240 ;
    END
  END l15_transducer_data_2[43]
  PIN l15_transducer_data_2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.490 2496.000 2157.770 2500.000 ;
    END
  END l15_transducer_data_2[44]
  PIN l15_transducer_data_2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 2496.000 2099.810 2500.000 ;
    END
  END l15_transducer_data_2[45]
  PIN l15_transducer_data_2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 785.440 2500.000 786.040 ;
    END
  END l15_transducer_data_2[46]
  PIN l15_transducer_data_2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 2496.000 1033.990 2500.000 ;
    END
  END l15_transducer_data_2[47]
  PIN l15_transducer_data_2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END l15_transducer_data_2[48]
  PIN l15_transducer_data_2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 2496.000 64.770 2500.000 ;
    END
  END l15_transducer_data_2[49]
  PIN l15_transducer_data_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 4.000 ;
    END
  END l15_transducer_data_2[4]
  PIN l15_transducer_data_2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END l15_transducer_data_2[50]
  PIN l15_transducer_data_2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END l15_transducer_data_2[51]
  PIN l15_transducer_data_2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END l15_transducer_data_2[52]
  PIN l15_transducer_data_2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 2496.000 1710.190 2500.000 ;
    END
  END l15_transducer_data_2[53]
  PIN l15_transducer_data_2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 884.040 2500.000 884.640 ;
    END
  END l15_transducer_data_2[54]
  PIN l15_transducer_data_2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 843.240 2500.000 843.840 ;
    END
  END l15_transducer_data_2[55]
  PIN l15_transducer_data_2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END l15_transducer_data_2[56]
  PIN l15_transducer_data_2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END l15_transducer_data_2[57]
  PIN l15_transducer_data_2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 2496.000 1307.690 2500.000 ;
    END
  END l15_transducer_data_2[58]
  PIN l15_transducer_data_2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END l15_transducer_data_2[59]
  PIN l15_transducer_data_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.390 0.000 2463.670 4.000 ;
    END
  END l15_transducer_data_2[5]
  PIN l15_transducer_data_2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 2496.000 1916.270 2500.000 ;
    END
  END l15_transducer_data_2[60]
  PIN l15_transducer_data_2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1519.840 2500.000 1520.440 ;
    END
  END l15_transducer_data_2[61]
  PIN l15_transducer_data_2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2461.640 4.000 2462.240 ;
    END
  END l15_transducer_data_2[62]
  PIN l15_transducer_data_2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2407.240 4.000 2407.840 ;
    END
  END l15_transducer_data_2[63]
  PIN l15_transducer_data_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 4.000 ;
    END
  END l15_transducer_data_2[6]
  PIN l15_transducer_data_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1938.040 4.000 1938.640 ;
    END
  END l15_transducer_data_2[7]
  PIN l15_transducer_data_2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END l15_transducer_data_2[8]
  PIN l15_transducer_data_2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.150 2496.000 2489.430 2500.000 ;
    END
  END l15_transducer_data_2[9]
  PIN l15_transducer_data_3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 2496.000 2012.870 2500.000 ;
    END
  END l15_transducer_data_3[0]
  PIN l15_transducer_data_3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1730.640 2500.000 1731.240 ;
    END
  END l15_transducer_data_3[10]
  PIN l15_transducer_data_3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 686.840 2500.000 687.440 ;
    END
  END l15_transducer_data_3[11]
  PIN l15_transducer_data_3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END l15_transducer_data_3[12]
  PIN l15_transducer_data_3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END l15_transducer_data_3[13]
  PIN l15_transducer_data_3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END l15_transducer_data_3[14]
  PIN l15_transducer_data_3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END l15_transducer_data_3[15]
  PIN l15_transducer_data_3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END l15_transducer_data_3[16]
  PIN l15_transducer_data_3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1067.640 2500.000 1068.240 ;
    END
  END l15_transducer_data_3[17]
  PIN l15_transducer_data_3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2417.440 2500.000 2418.040 ;
    END
  END l15_transducer_data_3[18]
  PIN l15_transducer_data_3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END l15_transducer_data_3[19]
  PIN l15_transducer_data_3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 0.000 1658.670 4.000 ;
    END
  END l15_transducer_data_3[1]
  PIN l15_transducer_data_3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.870 0.000 2090.150 4.000 ;
    END
  END l15_transducer_data_3[20]
  PIN l15_transducer_data_3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 2496.000 1439.710 2500.000 ;
    END
  END l15_transducer_data_3[21]
  PIN l15_transducer_data_3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END l15_transducer_data_3[22]
  PIN l15_transducer_data_3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.040 4.000 1530.640 ;
    END
  END l15_transducer_data_3[23]
  PIN l15_transducer_data_3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 17.040 2500.000 17.640 ;
    END
  END l15_transducer_data_3[24]
  PIN l15_transducer_data_3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END l15_transducer_data_3[25]
  PIN l15_transducer_data_3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1734.040 2500.000 1734.640 ;
    END
  END l15_transducer_data_3[26]
  PIN l15_transducer_data_3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 295.840 2500.000 296.440 ;
    END
  END l15_transducer_data_3[27]
  PIN l15_transducer_data_3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 4.000 1415.040 ;
    END
  END l15_transducer_data_3[28]
  PIN l15_transducer_data_3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 2496.000 1008.230 2500.000 ;
    END
  END l15_transducer_data_3[29]
  PIN l15_transducer_data_3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END l15_transducer_data_3[2]
  PIN l15_transducer_data_3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END l15_transducer_data_3[30]
  PIN l15_transducer_data_3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 0.000 1935.590 4.000 ;
    END
  END l15_transducer_data_3[31]
  PIN l15_transducer_data_3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END l15_transducer_data_3[32]
  PIN l15_transducer_data_3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 2496.000 702.330 2500.000 ;
    END
  END l15_transducer_data_3[33]
  PIN l15_transducer_data_3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2196.440 2500.000 2197.040 ;
    END
  END l15_transducer_data_3[34]
  PIN l15_transducer_data_3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 2496.000 863.330 2500.000 ;
    END
  END l15_transducer_data_3[35]
  PIN l15_transducer_data_3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.890 0.000 2222.170 4.000 ;
    END
  END l15_transducer_data_3[36]
  PIN l15_transducer_data_3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2237.240 4.000 2237.840 ;
    END
  END l15_transducer_data_3[37]
  PIN l15_transducer_data_3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1808.840 2500.000 1809.440 ;
    END
  END l15_transducer_data_3[38]
  PIN l15_transducer_data_3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END l15_transducer_data_3[39]
  PIN l15_transducer_data_3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1179.840 2500.000 1180.440 ;
    END
  END l15_transducer_data_3[3]
  PIN l15_transducer_data_3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 51.040 2500.000 51.640 ;
    END
  END l15_transducer_data_3[40]
  PIN l15_transducer_data_3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END l15_transducer_data_3[41]
  PIN l15_transducer_data_3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END l15_transducer_data_3[42]
  PIN l15_transducer_data_3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2111.440 2500.000 2112.040 ;
    END
  END l15_transducer_data_3[43]
  PIN l15_transducer_data_3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 962.240 2500.000 962.840 ;
    END
  END l15_transducer_data_3[44]
  PIN l15_transducer_data_3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END l15_transducer_data_3[45]
  PIN l15_transducer_data_3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2125.040 2500.000 2125.640 ;
    END
  END l15_transducer_data_3[46]
  PIN l15_transducer_data_3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END l15_transducer_data_3[47]
  PIN l15_transducer_data_3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END l15_transducer_data_3[48]
  PIN l15_transducer_data_3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 142.840 2500.000 143.440 ;
    END
  END l15_transducer_data_3[49]
  PIN l15_transducer_data_3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END l15_transducer_data_3[4]
  PIN l15_transducer_data_3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 2496.000 415.750 2500.000 ;
    END
  END l15_transducer_data_3[50]
  PIN l15_transducer_data_3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END l15_transducer_data_3[51]
  PIN l15_transducer_data_3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 2496.000 1146.690 2500.000 ;
    END
  END l15_transducer_data_3[52]
  PIN l15_transducer_data_3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 635.840 2500.000 636.440 ;
    END
  END l15_transducer_data_3[53]
  PIN l15_transducer_data_3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 2496.000 1874.410 2500.000 ;
    END
  END l15_transducer_data_3[54]
  PIN l15_transducer_data_3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END l15_transducer_data_3[55]
  PIN l15_transducer_data_3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.630 2496.000 2276.910 2500.000 ;
    END
  END l15_transducer_data_3[56]
  PIN l15_transducer_data_3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END l15_transducer_data_3[57]
  PIN l15_transducer_data_3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 2496.000 1108.050 2500.000 ;
    END
  END l15_transducer_data_3[58]
  PIN l15_transducer_data_3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.070 2496.000 2444.350 2500.000 ;
    END
  END l15_transducer_data_3[59]
  PIN l15_transducer_data_3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1513.040 2500.000 1513.640 ;
    END
  END l15_transducer_data_3[5]
  PIN l15_transducer_data_3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END l15_transducer_data_3[60]
  PIN l15_transducer_data_3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1598.040 2500.000 1598.640 ;
    END
  END l15_transducer_data_3[61]
  PIN l15_transducer_data_3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END l15_transducer_data_3[62]
  PIN l15_transducer_data_3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 2496.000 187.130 2500.000 ;
    END
  END l15_transducer_data_3[63]
  PIN l15_transducer_data_3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2434.440 2500.000 2435.040 ;
    END
  END l15_transducer_data_3[6]
  PIN l15_transducer_data_3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 2496.000 544.550 2500.000 ;
    END
  END l15_transducer_data_3[7]
  PIN l15_transducer_data_3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1907.440 4.000 1908.040 ;
    END
  END l15_transducer_data_3[8]
  PIN l15_transducer_data_3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END l15_transducer_data_3[9]
  PIN l15_transducer_error[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 850.040 2500.000 850.640 ;
    END
  END l15_transducer_error[0]
  PIN l15_transducer_error[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 2496.000 988.910 2500.000 ;
    END
  END l15_transducer_error[1]
  PIN l15_transducer_f4b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.240 4.000 1914.840 ;
    END
  END l15_transducer_f4b
  PIN l15_transducer_header_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 4.000 ;
    END
  END l15_transducer_header_ack
  PIN l15_transducer_inval_address_15_4[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1965.240 2500.000 1965.840 ;
    END
  END l15_transducer_inval_address_15_4[10]
  PIN l15_transducer_inval_address_15_4[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 353.640 2500.000 354.240 ;
    END
  END l15_transducer_inval_address_15_4[11]
  PIN l15_transducer_inval_address_15_4[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END l15_transducer_inval_address_15_4[12]
  PIN l15_transducer_inval_address_15_4[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 2496.000 1816.450 2500.000 ;
    END
  END l15_transducer_inval_address_15_4[13]
  PIN l15_transducer_inval_address_15_4[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END l15_transducer_inval_address_15_4[14]
  PIN l15_transducer_inval_address_15_4[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END l15_transducer_inval_address_15_4[15]
  PIN l15_transducer_inval_address_15_4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 2496.000 650.810 2500.000 ;
    END
  END l15_transducer_inval_address_15_4[4]
  PIN l15_transducer_inval_address_15_4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 2496.000 1504.110 2500.000 ;
    END
  END l15_transducer_inval_address_15_4[5]
  PIN l15_transducer_inval_address_15_4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 54.440 2500.000 55.040 ;
    END
  END l15_transducer_inval_address_15_4[6]
  PIN l15_transducer_inval_address_15_4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 2496.000 418.970 2500.000 ;
    END
  END l15_transducer_inval_address_15_4[7]
  PIN l15_transducer_inval_address_15_4[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.810 0.000 2338.090 4.000 ;
    END
  END l15_transducer_inval_address_15_4[8]
  PIN l15_transducer_inval_address_15_4[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1700.040 2500.000 1700.640 ;
    END
  END l15_transducer_inval_address_15_4[9]
  PIN l15_transducer_inval_dcache_all_way
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 4.000 ;
    END
  END l15_transducer_inval_dcache_all_way
  PIN l15_transducer_inval_dcache_inval
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END l15_transducer_inval_dcache_inval
  PIN l15_transducer_inval_icache_all_way
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END l15_transducer_inval_icache_all_way
  PIN l15_transducer_inval_icache_inval
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1978.840 4.000 1979.440 ;
    END
  END l15_transducer_inval_icache_inval
  PIN l15_transducer_inval_way[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END l15_transducer_inval_way[0]
  PIN l15_transducer_inval_way[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.490 2496.000 2479.770 2500.000 ;
    END
  END l15_transducer_inval_way[1]
  PIN l15_transducer_l2miss
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END l15_transducer_l2miss
  PIN l15_transducer_noncacheable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END l15_transducer_noncacheable
  PIN l15_transducer_prefetch
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END l15_transducer_prefetch
  PIN l15_transducer_returntype[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2152.240 2500.000 2152.840 ;
    END
  END l15_transducer_returntype[0]
  PIN l15_transducer_returntype[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2458.240 4.000 2458.840 ;
    END
  END l15_transducer_returntype[1]
  PIN l15_transducer_returntype[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.390 2496.000 1819.670 2500.000 ;
    END
  END l15_transducer_returntype[2]
  PIN l15_transducer_returntype[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 2496.000 634.710 2500.000 ;
    END
  END l15_transducer_returntype[3]
  PIN l15_transducer_threadid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2397.040 4.000 2397.640 ;
    END
  END l15_transducer_threadid
  PIN l15_transducer_val
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 683.440 2500.000 684.040 ;
    END
  END l15_transducer_val
  PIN l2_rtap_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END l2_rtap_data[0]
  PIN l2_rtap_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END l2_rtap_data[1]
  PIN l2_rtap_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END l2_rtap_data[2]
  PIN l2_rtap_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1455.240 2500.000 1455.840 ;
    END
  END l2_rtap_data[3]
  PIN noc1_out_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END noc1_out_data[0]
  PIN noc1_out_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END noc1_out_data[10]
  PIN noc1_out_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 2496.000 557.430 2500.000 ;
    END
  END noc1_out_data[11]
  PIN noc1_out_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END noc1_out_data[12]
  PIN noc1_out_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 615.440 2500.000 616.040 ;
    END
  END noc1_out_data[13]
  PIN noc1_out_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.290 0.000 2447.570 4.000 ;
    END
  END noc1_out_data[14]
  PIN noc1_out_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.350 0.000 2360.630 4.000 ;
    END
  END noc1_out_data[15]
  PIN noc1_out_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END noc1_out_data[16]
  PIN noc1_out_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 2496.000 522.010 2500.000 ;
    END
  END noc1_out_data[17]
  PIN noc1_out_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1972.040 4.000 1972.640 ;
    END
  END noc1_out_data[18]
  PIN noc1_out_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2108.040 4.000 2108.640 ;
    END
  END noc1_out_data[19]
  PIN noc1_out_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2213.440 2500.000 2214.040 ;
    END
  END noc1_out_data[1]
  PIN noc1_out_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2077.440 4.000 2078.040 ;
    END
  END noc1_out_data[20]
  PIN noc1_out_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2053.640 2500.000 2054.240 ;
    END
  END noc1_out_data[21]
  PIN noc1_out_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 996.240 2500.000 996.840 ;
    END
  END noc1_out_data[22]
  PIN noc1_out_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 166.640 2500.000 167.240 ;
    END
  END noc1_out_data[23]
  PIN noc1_out_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2390.240 4.000 2390.840 ;
    END
  END noc1_out_data[24]
  PIN noc1_out_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END noc1_out_data[25]
  PIN noc1_out_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END noc1_out_data[26]
  PIN noc1_out_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 2496.000 1339.890 2500.000 ;
    END
  END noc1_out_data[27]
  PIN noc1_out_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 510.040 2500.000 510.640 ;
    END
  END noc1_out_data[28]
  PIN noc1_out_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 2496.000 235.430 2500.000 ;
    END
  END noc1_out_data[29]
  PIN noc1_out_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2482.040 4.000 2482.640 ;
    END
  END noc1_out_data[2]
  PIN noc1_out_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 0.000 2257.590 4.000 ;
    END
  END noc1_out_data[30]
  PIN noc1_out_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2142.040 4.000 2142.640 ;
    END
  END noc1_out_data[31]
  PIN noc1_out_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1370.240 2500.000 1370.840 ;
    END
  END noc1_out_data[32]
  PIN noc1_out_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2250.840 4.000 2251.440 ;
    END
  END noc1_out_data[33]
  PIN noc1_out_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1781.640 4.000 1782.240 ;
    END
  END noc1_out_data[34]
  PIN noc1_out_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END noc1_out_data[35]
  PIN noc1_out_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END noc1_out_data[36]
  PIN noc1_out_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 2496.000 2138.450 2500.000 ;
    END
  END noc1_out_data[37]
  PIN noc1_out_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 2496.000 1140.250 2500.000 ;
    END
  END noc1_out_data[38]
  PIN noc1_out_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END noc1_out_data[39]
  PIN noc1_out_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2257.640 2500.000 2258.240 ;
    END
  END noc1_out_data[3]
  PIN noc1_out_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.630 0.000 2276.910 4.000 ;
    END
  END noc1_out_data[40]
  PIN noc1_out_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1638.840 2500.000 1639.440 ;
    END
  END noc1_out_data[41]
  PIN noc1_out_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 2496.000 1500.890 2500.000 ;
    END
  END noc1_out_data[42]
  PIN noc1_out_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END noc1_out_data[43]
  PIN noc1_out_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.240 4.000 1404.840 ;
    END
  END noc1_out_data[44]
  PIN noc1_out_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 2496.000 338.470 2500.000 ;
    END
  END noc1_out_data[45]
  PIN noc1_out_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1591.240 2500.000 1591.840 ;
    END
  END noc1_out_data[46]
  PIN noc1_out_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END noc1_out_data[47]
  PIN noc1_out_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2318.840 2500.000 2319.440 ;
    END
  END noc1_out_data[48]
  PIN noc1_out_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 2496.000 2115.910 2500.000 ;
    END
  END noc1_out_data[49]
  PIN noc1_out_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1683.040 2500.000 1683.640 ;
    END
  END noc1_out_data[4]
  PIN noc1_out_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 370.640 2500.000 371.240 ;
    END
  END noc1_out_data[50]
  PIN noc1_out_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END noc1_out_data[51]
  PIN noc1_out_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1101.640 2500.000 1102.240 ;
    END
  END noc1_out_data[52]
  PIN noc1_out_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 2496.000 2218.950 2500.000 ;
    END
  END noc1_out_data[53]
  PIN noc1_out_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2468.440 4.000 2469.040 ;
    END
  END noc1_out_data[54]
  PIN noc1_out_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 2496.000 77.650 2500.000 ;
    END
  END noc1_out_data[55]
  PIN noc1_out_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1557.240 2500.000 1557.840 ;
    END
  END noc1_out_data[56]
  PIN noc1_out_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 751.440 2500.000 752.040 ;
    END
  END noc1_out_data[57]
  PIN noc1_out_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1825.840 4.000 1826.440 ;
    END
  END noc1_out_data[58]
  PIN noc1_out_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1873.440 4.000 1874.040 ;
    END
  END noc1_out_data[59]
  PIN noc1_out_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2458.240 2500.000 2458.840 ;
    END
  END noc1_out_data[5]
  PIN noc1_out_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.490 0.000 1996.770 4.000 ;
    END
  END noc1_out_data[60]
  PIN noc1_out_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 0.000 2048.290 4.000 ;
    END
  END noc1_out_data[61]
  PIN noc1_out_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.590 0.000 2173.870 4.000 ;
    END
  END noc1_out_data[62]
  PIN noc1_out_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.050 2496.000 2151.330 2500.000 ;
    END
  END noc1_out_data[63]
  PIN noc1_out_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 540.640 2500.000 541.240 ;
    END
  END noc1_out_data[6]
  PIN noc1_out_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1768.040 2500.000 1768.640 ;
    END
  END noc1_out_data[7]
  PIN noc1_out_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END noc1_out_data[8]
  PIN noc1_out_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2063.840 2500.000 2064.440 ;
    END
  END noc1_out_data[9]
  PIN noc1_out_rdy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2291.640 2500.000 2292.240 ;
    END
  END noc1_out_rdy
  PIN noc1_out_val
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 30.640 2500.000 31.240 ;
    END
  END noc1_out_val
  PIN noc2_in_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 2496.000 1961.350 2500.000 ;
    END
  END noc2_in_data[0]
  PIN noc2_in_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 2496.000 1436.490 2500.000 ;
    END
  END noc2_in_data[10]
  PIN noc2_in_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 2496.000 377.110 2500.000 ;
    END
  END noc2_in_data[11]
  PIN noc2_in_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.790 2496.000 1240.070 2500.000 ;
    END
  END noc2_in_data[12]
  PIN noc2_in_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.810 2496.000 2016.090 2500.000 ;
    END
  END noc2_in_data[13]
  PIN noc2_in_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 544.040 2500.000 544.640 ;
    END
  END noc2_in_data[14]
  PIN noc2_in_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 2496.000 1211.090 2500.000 ;
    END
  END noc2_in_data[15]
  PIN noc2_in_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 4.000 ;
    END
  END noc2_in_data[16]
  PIN noc2_in_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 193.840 2500.000 194.440 ;
    END
  END noc2_in_data[17]
  PIN noc2_in_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1662.640 2500.000 1663.240 ;
    END
  END noc2_in_data[18]
  PIN noc2_in_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 0.000 1958.130 4.000 ;
    END
  END noc2_in_data[19]
  PIN noc2_in_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END noc2_in_data[1]
  PIN noc2_in_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END noc2_in_data[20]
  PIN noc2_in_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END noc2_in_data[21]
  PIN noc2_in_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END noc2_in_data[22]
  PIN noc2_in_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1591.240 4.000 1591.840 ;
    END
  END noc2_in_data[23]
  PIN noc2_in_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.730 2496.000 1971.010 2500.000 ;
    END
  END noc2_in_data[24]
  PIN noc2_in_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1281.840 2500.000 1282.440 ;
    END
  END noc2_in_data[25]
  PIN noc2_in_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 2496.000 1636.130 2500.000 ;
    END
  END noc2_in_data[26]
  PIN noc2_in_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1608.240 2500.000 1608.840 ;
    END
  END noc2_in_data[27]
  PIN noc2_in_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2162.440 2500.000 2163.040 ;
    END
  END noc2_in_data[28]
  PIN noc2_in_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 34.040 2500.000 34.640 ;
    END
  END noc2_in_data[29]
  PIN noc2_in_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END noc2_in_data[2]
  PIN noc2_in_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 0.000 2354.190 4.000 ;
    END
  END noc2_in_data[30]
  PIN noc2_in_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END noc2_in_data[31]
  PIN noc2_in_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1737.440 4.000 1738.040 ;
    END
  END noc2_in_data[32]
  PIN noc2_in_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 2496.000 1851.870 2500.000 ;
    END
  END noc2_in_data[33]
  PIN noc2_in_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2026.440 4.000 2027.040 ;
    END
  END noc2_in_data[34]
  PIN noc2_in_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END noc2_in_data[35]
  PIN noc2_in_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 629.040 2500.000 629.640 ;
    END
  END noc2_in_data[36]
  PIN noc2_in_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END noc2_in_data[37]
  PIN noc2_in_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2468.440 2500.000 2469.040 ;
    END
  END noc2_in_data[38]
  PIN noc2_in_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.270 2496.000 2315.550 2500.000 ;
    END
  END noc2_in_data[39]
  PIN noc2_in_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 2496.000 1793.910 2500.000 ;
    END
  END noc2_in_data[3]
  PIN noc2_in_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2366.440 4.000 2367.040 ;
    END
  END noc2_in_data[40]
  PIN noc2_in_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 2496.000 815.030 2500.000 ;
    END
  END noc2_in_data[41]
  PIN noc2_in_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END noc2_in_data[42]
  PIN noc2_in_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2029.840 4.000 2030.440 ;
    END
  END noc2_in_data[43]
  PIN noc2_in_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END noc2_in_data[44]
  PIN noc2_in_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 2496.000 254.750 2500.000 ;
    END
  END noc2_in_data[45]
  PIN noc2_in_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.930 2496.000 2003.210 2500.000 ;
    END
  END noc2_in_data[46]
  PIN noc2_in_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1397.440 4.000 1398.040 ;
    END
  END noc2_in_data[47]
  PIN noc2_in_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 2496.000 840.790 2500.000 ;
    END
  END noc2_in_data[48]
  PIN noc2_in_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 935.040 2500.000 935.640 ;
    END
  END noc2_in_data[49]
  PIN noc2_in_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2437.840 4.000 2438.440 ;
    END
  END noc2_in_data[4]
  PIN noc2_in_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 2496.000 190.350 2500.000 ;
    END
  END noc2_in_data[50]
  PIN noc2_in_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2342.640 4.000 2343.240 ;
    END
  END noc2_in_data[51]
  PIN noc2_in_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 2496.000 267.630 2500.000 ;
    END
  END noc2_in_data[52]
  PIN noc2_in_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END noc2_in_data[53]
  PIN noc2_in_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 2496.000 1491.230 2500.000 ;
    END
  END noc2_in_data[54]
  PIN noc2_in_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 455.640 2500.000 456.240 ;
    END
  END noc2_in_data[55]
  PIN noc2_in_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.030 0.000 2341.310 4.000 ;
    END
  END noc2_in_data[56]
  PIN noc2_in_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END noc2_in_data[57]
  PIN noc2_in_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END noc2_in_data[58]
  PIN noc2_in_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.790 2496.000 2045.070 2500.000 ;
    END
  END noc2_in_data[59]
  PIN noc2_in_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2441.240 4.000 2441.840 ;
    END
  END noc2_in_data[5]
  PIN noc2_in_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END noc2_in_data[60]
  PIN noc2_in_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2322.240 2500.000 2322.840 ;
    END
  END noc2_in_data[61]
  PIN noc2_in_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2301.840 4.000 2302.440 ;
    END
  END noc2_in_data[62]
  PIN noc2_in_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1689.840 4.000 1690.440 ;
    END
  END noc2_in_data[63]
  PIN noc2_in_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END noc2_in_data[6]
  PIN noc2_in_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END noc2_in_data[7]
  PIN noc2_in_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.350 0.000 2038.630 4.000 ;
    END
  END noc2_in_data[8]
  PIN noc2_in_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 0.000 2199.630 4.000 ;
    END
  END noc2_in_data[9]
  PIN noc2_in_rdy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2080.840 2500.000 2081.440 ;
    END
  END noc2_in_rdy
  PIN noc2_in_val
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END noc2_in_val
  PIN noc3_out_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2312.040 2500.000 2312.640 ;
    END
  END noc3_out_data[0]
  PIN noc3_out_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END noc3_out_data[10]
  PIN noc3_out_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 2496.000 457.610 2500.000 ;
    END
  END noc3_out_data[11]
  PIN noc3_out_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 0.000 1478.350 4.000 ;
    END
  END noc3_out_data[12]
  PIN noc3_out_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.750 2496.000 1781.030 2500.000 ;
    END
  END noc3_out_data[13]
  PIN noc3_out_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END noc3_out_data[14]
  PIN noc3_out_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 0.000 2183.530 4.000 ;
    END
  END noc3_out_data[15]
  PIN noc3_out_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 2496.000 1471.910 2500.000 ;
    END
  END noc3_out_data[16]
  PIN noc3_out_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END noc3_out_data[17]
  PIN noc3_out_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END noc3_out_data[18]
  PIN noc3_out_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1995.840 4.000 1996.440 ;
    END
  END noc3_out_data[19]
  PIN noc3_out_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.310 0.000 1774.590 4.000 ;
    END
  END noc3_out_data[1]
  PIN noc3_out_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END noc3_out_data[20]
  PIN noc3_out_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END noc3_out_data[21]
  PIN noc3_out_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 418.240 2500.000 418.840 ;
    END
  END noc3_out_data[22]
  PIN noc3_out_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 2496.000 1623.250 2500.000 ;
    END
  END noc3_out_data[23]
  PIN noc3_out_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END noc3_out_data[24]
  PIN noc3_out_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 2496.000 238.650 2500.000 ;
    END
  END noc3_out_data[25]
  PIN noc3_out_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1859.840 4.000 1860.440 ;
    END
  END noc3_out_data[26]
  PIN noc3_out_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2016.240 2500.000 2016.840 ;
    END
  END noc3_out_data[27]
  PIN noc3_out_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 836.440 2500.000 837.040 ;
    END
  END noc3_out_data[28]
  PIN noc3_out_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 938.440 2500.000 939.040 ;
    END
  END noc3_out_data[29]
  PIN noc3_out_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 2496.000 1478.350 2500.000 ;
    END
  END noc3_out_data[2]
  PIN noc3_out_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END noc3_out_data[30]
  PIN noc3_out_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 4.000 ;
    END
  END noc3_out_data[31]
  PIN noc3_out_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END noc3_out_data[32]
  PIN noc3_out_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 2496.000 1858.310 2500.000 ;
    END
  END noc3_out_data[33]
  PIN noc3_out_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END noc3_out_data[34]
  PIN noc3_out_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END noc3_out_data[35]
  PIN noc3_out_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 2496.000 444.730 2500.000 ;
    END
  END noc3_out_data[36]
  PIN noc3_out_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1985.640 2500.000 1986.240 ;
    END
  END noc3_out_data[37]
  PIN noc3_out_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 2496.000 1285.150 2500.000 ;
    END
  END noc3_out_data[38]
  PIN noc3_out_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END noc3_out_data[39]
  PIN noc3_out_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 4.000 ;
    END
  END noc3_out_data[3]
  PIN noc3_out_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 2496.000 1562.070 2500.000 ;
    END
  END noc3_out_data[40]
  PIN noc3_out_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 306.040 2500.000 306.640 ;
    END
  END noc3_out_data[41]
  PIN noc3_out_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.390 2496.000 2302.670 2500.000 ;
    END
  END noc3_out_data[42]
  PIN noc3_out_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 2496.000 3.590 2500.000 ;
    END
  END noc3_out_data[43]
  PIN noc3_out_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END noc3_out_data[44]
  PIN noc3_out_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 2496.000 1394.630 2500.000 ;
    END
  END noc3_out_data[45]
  PIN noc3_out_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 4.000 ;
    END
  END noc3_out_data[46]
  PIN noc3_out_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1972.040 2500.000 1972.640 ;
    END
  END noc3_out_data[47]
  PIN noc3_out_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 268.640 2500.000 269.240 ;
    END
  END noc3_out_data[48]
  PIN noc3_out_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END noc3_out_data[49]
  PIN noc3_out_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 2496.000 180.690 2500.000 ;
    END
  END noc3_out_data[4]
  PIN noc3_out_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 2496.000 496.250 2500.000 ;
    END
  END noc3_out_data[50]
  PIN noc3_out_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END noc3_out_data[51]
  PIN noc3_out_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 2496.000 335.250 2500.000 ;
    END
  END noc3_out_data[52]
  PIN noc3_out_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2233.840 2500.000 2234.440 ;
    END
  END noc3_out_data[53]
  PIN noc3_out_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 989.440 2500.000 990.040 ;
    END
  END noc3_out_data[54]
  PIN noc3_out_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.330 2496.000 1906.610 2500.000 ;
    END
  END noc3_out_data[55]
  PIN noc3_out_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1322.640 4.000 1323.240 ;
    END
  END noc3_out_data[56]
  PIN noc3_out_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 2496.000 1913.050 2500.000 ;
    END
  END noc3_out_data[57]
  PIN noc3_out_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1645.640 2500.000 1646.240 ;
    END
  END noc3_out_data[58]
  PIN noc3_out_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 710.640 2500.000 711.240 ;
    END
  END noc3_out_data[59]
  PIN noc3_out_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 2496.000 428.630 2500.000 ;
    END
  END noc3_out_data[5]
  PIN noc3_out_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END noc3_out_data[60]
  PIN noc3_out_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.090 0.000 2093.370 4.000 ;
    END
  END noc3_out_data[61]
  PIN noc3_out_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.450 0.000 2054.730 4.000 ;
    END
  END noc3_out_data[62]
  PIN noc3_out_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 734.440 2500.000 735.040 ;
    END
  END noc3_out_data[63]
  PIN noc3_out_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 2496.000 776.390 2500.000 ;
    END
  END noc3_out_data[6]
  PIN noc3_out_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END noc3_out_data[7]
  PIN noc3_out_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 2496.000 1545.970 2500.000 ;
    END
  END noc3_out_data[8]
  PIN noc3_out_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.550 2496.000 2231.830 2500.000 ;
    END
  END noc3_out_data[9]
  PIN noc3_out_rdy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.310 0.000 2096.590 4.000 ;
    END
  END noc3_out_rdy
  PIN noc3_out_val
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2424.240 2500.000 2424.840 ;
    END
  END noc3_out_val
  PIN processor_router_data_noc2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.240 4.000 1251.840 ;
    END
  END processor_router_data_noc2[0]
  PIN processor_router_data_noc2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1462.040 2500.000 1462.640 ;
    END
  END processor_router_data_noc2[10]
  PIN processor_router_data_noc2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1846.240 2500.000 1846.840 ;
    END
  END processor_router_data_noc2[11]
  PIN processor_router_data_noc2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2227.040 2500.000 2227.640 ;
    END
  END processor_router_data_noc2[12]
  PIN processor_router_data_noc2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END processor_router_data_noc2[13]
  PIN processor_router_data_noc2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 2496.000 1449.370 2500.000 ;
    END
  END processor_router_data_noc2[14]
  PIN processor_router_data_noc2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.430 0.000 2083.710 4.000 ;
    END
  END processor_router_data_noc2[15]
  PIN processor_router_data_noc2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 2496.000 1848.650 2500.000 ;
    END
  END processor_router_data_noc2[16]
  PIN processor_router_data_noc2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END processor_router_data_noc2[17]
  PIN processor_router_data_noc2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 530.440 2500.000 531.040 ;
    END
  END processor_router_data_noc2[18]
  PIN processor_router_data_noc2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.970 0.000 2428.250 4.000 ;
    END
  END processor_router_data_noc2[19]
  PIN processor_router_data_noc2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END processor_router_data_noc2[1]
  PIN processor_router_data_noc2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END processor_router_data_noc2[20]
  PIN processor_router_data_noc2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1142.440 2500.000 1143.040 ;
    END
  END processor_router_data_noc2[21]
  PIN processor_router_data_noc2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1989.040 2500.000 1989.640 ;
    END
  END processor_router_data_noc2[22]
  PIN processor_router_data_noc2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END processor_router_data_noc2[23]
  PIN processor_router_data_noc2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 2496.000 2048.290 2500.000 ;
    END
  END processor_router_data_noc2[24]
  PIN processor_router_data_noc2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 0.000 2328.430 4.000 ;
    END
  END processor_router_data_noc2[25]
  PIN processor_router_data_noc2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END processor_router_data_noc2[26]
  PIN processor_router_data_noc2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END processor_router_data_noc2[27]
  PIN processor_router_data_noc2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.150 0.000 2489.430 4.000 ;
    END
  END processor_router_data_noc2[28]
  PIN processor_router_data_noc2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END processor_router_data_noc2[29]
  PIN processor_router_data_noc2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 139.440 2500.000 140.040 ;
    END
  END processor_router_data_noc2[2]
  PIN processor_router_data_noc2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 2496.000 1130.590 2500.000 ;
    END
  END processor_router_data_noc2[30]
  PIN processor_router_data_noc2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1955.040 2500.000 1955.640 ;
    END
  END processor_router_data_noc2[31]
  PIN processor_router_data_noc2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 2496.000 1265.830 2500.000 ;
    END
  END processor_router_data_noc2[32]
  PIN processor_router_data_noc2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.010 0.000 2209.290 4.000 ;
    END
  END processor_router_data_noc2[33]
  PIN processor_router_data_noc2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.930 0.000 2164.210 4.000 ;
    END
  END processor_router_data_noc2[34]
  PIN processor_router_data_noc2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END processor_router_data_noc2[35]
  PIN processor_router_data_noc2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END processor_router_data_noc2[36]
  PIN processor_router_data_noc2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1271.640 4.000 1272.240 ;
    END
  END processor_router_data_noc2[37]
  PIN processor_router_data_noc2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END processor_router_data_noc2[38]
  PIN processor_router_data_noc2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 731.040 2500.000 731.640 ;
    END
  END processor_router_data_noc2[39]
  PIN processor_router_data_noc2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1108.440 2500.000 1109.040 ;
    END
  END processor_router_data_noc2[3]
  PIN processor_router_data_noc2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 2496.000 1185.330 2500.000 ;
    END
  END processor_router_data_noc2[40]
  PIN processor_router_data_noc2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END processor_router_data_noc2[41]
  PIN processor_router_data_noc2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2182.840 2500.000 2183.440 ;
    END
  END processor_router_data_noc2[42]
  PIN processor_router_data_noc2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.650 0.000 1925.930 4.000 ;
    END
  END processor_router_data_noc2[43]
  PIN processor_router_data_noc2[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END processor_router_data_noc2[44]
  PIN processor_router_data_noc2[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 0.000 1481.570 4.000 ;
    END
  END processor_router_data_noc2[45]
  PIN processor_router_data_noc2[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END processor_router_data_noc2[46]
  PIN processor_router_data_noc2[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.270 0.000 2154.550 4.000 ;
    END
  END processor_router_data_noc2[47]
  PIN processor_router_data_noc2[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 503.240 2500.000 503.840 ;
    END
  END processor_router_data_noc2[48]
  PIN processor_router_data_noc2[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.450 0.000 2376.730 4.000 ;
    END
  END processor_router_data_noc2[49]
  PIN processor_router_data_noc2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END processor_router_data_noc2[4]
  PIN processor_router_data_noc2[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 2496.000 1252.950 2500.000 ;
    END
  END processor_router_data_noc2[50]
  PIN processor_router_data_noc2[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 0.000 1961.350 4.000 ;
    END
  END processor_router_data_noc2[51]
  PIN processor_router_data_noc2[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1883.640 2500.000 1884.240 ;
    END
  END processor_router_data_noc2[52]
  PIN processor_router_data_noc2[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END processor_router_data_noc2[53]
  PIN processor_router_data_noc2[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2349.440 2500.000 2350.040 ;
    END
  END processor_router_data_noc2[54]
  PIN processor_router_data_noc2[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2131.840 2500.000 2132.440 ;
    END
  END processor_router_data_noc2[55]
  PIN processor_router_data_noc2[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END processor_router_data_noc2[56]
  PIN processor_router_data_noc2[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END processor_router_data_noc2[57]
  PIN processor_router_data_noc2[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 207.440 2500.000 208.040 ;
    END
  END processor_router_data_noc2[58]
  PIN processor_router_data_noc2[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2227.040 4.000 2227.640 ;
    END
  END processor_router_data_noc2[59]
  PIN processor_router_data_noc2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 656.240 2500.000 656.840 ;
    END
  END processor_router_data_noc2[5]
  PIN processor_router_data_noc2[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 2496.000 113.070 2500.000 ;
    END
  END processor_router_data_noc2[60]
  PIN processor_router_data_noc2[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END processor_router_data_noc2[61]
  PIN processor_router_data_noc2[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1360.040 2500.000 1360.640 ;
    END
  END processor_router_data_noc2[62]
  PIN processor_router_data_noc2[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 2496.000 1616.810 2500.000 ;
    END
  END processor_router_data_noc2[63]
  PIN processor_router_data_noc2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.250 0.000 2022.530 4.000 ;
    END
  END processor_router_data_noc2[6]
  PIN processor_router_data_noc2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2418.310 0.000 2418.590 4.000 ;
    END
  END processor_router_data_noc2[7]
  PIN processor_router_data_noc2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END processor_router_data_noc2[8]
  PIN processor_router_data_noc2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1764.640 4.000 1765.240 ;
    END
  END processor_router_data_noc2[9]
  PIN processor_router_ready_noc1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 346.840 2500.000 347.440 ;
    END
  END processor_router_ready_noc1
  PIN processor_router_ready_noc3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 703.840 2500.000 704.440 ;
    END
  END processor_router_ready_noc3
  PIN processor_router_valid_noc2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1856.440 4.000 1857.040 ;
    END
  END processor_router_valid_noc2
  PIN router_processor_ready_noc2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END router_processor_ready_noc2
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 2496.000 171.030 2500.000 ;
    END
  END rst_n
  PIN rtap_srams_bist_command[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 411.440 2500.000 412.040 ;
    END
  END rtap_srams_bist_command[0]
  PIN rtap_srams_bist_command[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2437.840 2500.000 2438.440 ;
    END
  END rtap_srams_bist_command[1]
  PIN rtap_srams_bist_command[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1961.840 4.000 1962.440 ;
    END
  END rtap_srams_bist_command[2]
  PIN rtap_srams_bist_command[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1870.040 4.000 1870.640 ;
    END
  END rtap_srams_bist_command[3]
  PIN rtap_srams_bist_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1285.240 2500.000 1285.840 ;
    END
  END rtap_srams_bist_data[0]
  PIN rtap_srams_bist_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.830 0.000 1665.110 4.000 ;
    END
  END rtap_srams_bist_data[1]
  PIN rtap_srams_bist_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.410 0.000 1951.690 4.000 ;
    END
  END rtap_srams_bist_data[2]
  PIN rtap_srams_bist_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 2496.000 183.910 2500.000 ;
    END
  END rtap_srams_bist_data[3]
  PIN srams_rtap_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1669.440 2500.000 1670.040 ;
    END
  END srams_rtap_data[0]
  PIN srams_rtap_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2046.840 4.000 2047.440 ;
    END
  END srams_rtap_data[1]
  PIN srams_rtap_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END srams_rtap_data[2]
  PIN srams_rtap_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 2496.000 1700.530 2500.000 ;
    END
  END srams_rtap_data[3]
  PIN tile_jtag_ucb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 153.040 2500.000 153.640 ;
    END
  END tile_jtag_ucb_data[0]
  PIN tile_jtag_ucb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 2496.000 125.950 2500.000 ;
    END
  END tile_jtag_ucb_data[1]
  PIN tile_jtag_ucb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 2496.000 1771.370 2500.000 ;
    END
  END tile_jtag_ucb_data[2]
  PIN tile_jtag_ucb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END tile_jtag_ucb_data[3]
  PIN tile_jtag_ucb_val
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1941.440 4.000 1942.040 ;
    END
  END tile_jtag_ucb_val
  PIN transducer_l15_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END transducer_l15_address[0]
  PIN transducer_l15_address[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.530 2496.000 1133.810 2500.000 ;
    END
  END transducer_l15_address[10]
  PIN transducer_l15_address[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 102.040 2500.000 102.640 ;
    END
  END transducer_l15_address[11]
  PIN transducer_l15_address[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.050 2496.000 1990.330 2500.000 ;
    END
  END transducer_l15_address[12]
  PIN transducer_l15_address[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END transducer_l15_address[13]
  PIN transducer_l15_address[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END transducer_l15_address[14]
  PIN transducer_l15_address[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.670 0.000 2057.950 4.000 ;
    END
  END transducer_l15_address[15]
  PIN transducer_l15_address[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 4.000 ;
    END
  END transducer_l15_address[16]
  PIN transducer_l15_address[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 2496.000 567.090 2500.000 ;
    END
  END transducer_l15_address[17]
  PIN transducer_l15_address[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2492.240 2500.000 2492.840 ;
    END
  END transducer_l15_address[18]
  PIN transducer_l15_address[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1261.440 2500.000 1262.040 ;
    END
  END transducer_l15_address[19]
  PIN transducer_l15_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 2496.000 1922.710 2500.000 ;
    END
  END transducer_l15_address[1]
  PIN transducer_l15_address[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.430 0.000 2244.710 4.000 ;
    END
  END transducer_l15_address[20]
  PIN transducer_l15_address[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END transducer_l15_address[21]
  PIN transducer_l15_address[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1635.440 4.000 1636.040 ;
    END
  END transducer_l15_address[22]
  PIN transducer_l15_address[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 2496.000 1091.950 2500.000 ;
    END
  END transducer_l15_address[23]
  PIN transducer_l15_address[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2206.640 2500.000 2207.240 ;
    END
  END transducer_l15_address[24]
  PIN transducer_l15_address[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.070 2496.000 2283.350 2500.000 ;
    END
  END transducer_l15_address[25]
  PIN transducer_l15_address[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 357.040 2500.000 357.640 ;
    END
  END transducer_l15_address[26]
  PIN transducer_l15_address[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1893.840 2500.000 1894.440 ;
    END
  END transducer_l15_address[27]
  PIN transducer_l15_address[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 2496.000 1613.590 2500.000 ;
    END
  END transducer_l15_address[28]
  PIN transducer_l15_address[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.840 4.000 1724.440 ;
    END
  END transducer_l15_address[29]
  PIN transducer_l15_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END transducer_l15_address[2]
  PIN transducer_l15_address[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 0.000 1822.890 4.000 ;
    END
  END transducer_l15_address[30]
  PIN transducer_l15_address[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END transducer_l15_address[31]
  PIN transducer_l15_address[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1560.640 2500.000 1561.240 ;
    END
  END transducer_l15_address[32]
  PIN transducer_l15_address[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END transducer_l15_address[33]
  PIN transducer_l15_address[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END transducer_l15_address[34]
  PIN transducer_l15_address[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1451.840 2500.000 1452.440 ;
    END
  END transducer_l15_address[35]
  PIN transducer_l15_address[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 2496.000 921.290 2500.000 ;
    END
  END transducer_l15_address[36]
  PIN transducer_l15_address[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2369.840 2500.000 2370.440 ;
    END
  END transducer_l15_address[37]
  PIN transducer_l15_address[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END transducer_l15_address[38]
  PIN transducer_l15_address[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2094.440 2500.000 2095.040 ;
    END
  END transducer_l15_address[39]
  PIN transducer_l15_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.930 0.000 2325.210 4.000 ;
    END
  END transducer_l15_address[3]
  PIN transducer_l15_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 2496.000 361.010 2500.000 ;
    END
  END transducer_l15_address[4]
  PIN transducer_l15_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.610 0.000 2144.890 4.000 ;
    END
  END transducer_l15_address[5]
  PIN transducer_l15_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.750 2496.000 2264.030 2500.000 ;
    END
  END transducer_l15_address[6]
  PIN transducer_l15_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 2496.000 798.930 2500.000 ;
    END
  END transducer_l15_address[7]
  PIN transducer_l15_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 2496.000 441.510 2500.000 ;
    END
  END transducer_l15_address[8]
  PIN transducer_l15_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 4.000 2118.840 ;
    END
  END transducer_l15_address[9]
  PIN transducer_l15_amo_op[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 2496.000 872.990 2500.000 ;
    END
  END transducer_l15_amo_op[0]
  PIN transducer_l15_amo_op[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END transducer_l15_amo_op[1]
  PIN transducer_l15_amo_op[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END transducer_l15_amo_op[2]
  PIN transducer_l15_amo_op[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1047.240 2500.000 1047.840 ;
    END
  END transducer_l15_amo_op[3]
  PIN transducer_l15_blockinitstore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1910.840 2500.000 1911.440 ;
    END
  END transducer_l15_blockinitstore
  PIN transducer_l15_blockstore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 2496.000 2247.930 2500.000 ;
    END
  END transducer_l15_blockstore
  PIN transducer_l15_csm_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END transducer_l15_csm_data[0]
  PIN transducer_l15_csm_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 6.840 2500.000 7.440 ;
    END
  END transducer_l15_csm_data[10]
  PIN transducer_l15_csm_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 2496.000 1542.750 2500.000 ;
    END
  END transducer_l15_csm_data[11]
  PIN transducer_l15_csm_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.290 2496.000 1964.570 2500.000 ;
    END
  END transducer_l15_csm_data[12]
  PIN transducer_l15_csm_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 2496.000 695.890 2500.000 ;
    END
  END transducer_l15_csm_data[13]
  PIN transducer_l15_csm_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 2496.000 1278.710 2500.000 ;
    END
  END transducer_l15_csm_data[14]
  PIN transducer_l15_csm_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 499.840 2500.000 500.440 ;
    END
  END transducer_l15_csm_data[15]
  PIN transducer_l15_csm_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 2496.000 1246.510 2500.000 ;
    END
  END transducer_l15_csm_data[16]
  PIN transducer_l15_csm_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 363.840 2500.000 364.440 ;
    END
  END transducer_l15_csm_data[17]
  PIN transducer_l15_csm_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 945.240 2500.000 945.840 ;
    END
  END transducer_l15_csm_data[18]
  PIN transducer_l15_csm_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END transducer_l15_csm_data[19]
  PIN transducer_l15_csm_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END transducer_l15_csm_data[1]
  PIN transducer_l15_csm_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END transducer_l15_csm_data[20]
  PIN transducer_l15_csm_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1713.640 2500.000 1714.240 ;
    END
  END transducer_l15_csm_data[21]
  PIN transducer_l15_csm_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 2496.000 1649.010 2500.000 ;
    END
  END transducer_l15_csm_data[22]
  PIN transducer_l15_csm_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2040.040 4.000 2040.640 ;
    END
  END transducer_l15_csm_data[23]
  PIN transducer_l15_csm_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1910.840 4.000 1911.440 ;
    END
  END transducer_l15_csm_data[24]
  PIN transducer_l15_csm_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END transducer_l15_csm_data[25]
  PIN transducer_l15_csm_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END transducer_l15_csm_data[26]
  PIN transducer_l15_csm_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 2496.000 1381.750 2500.000 ;
    END
  END transducer_l15_csm_data[27]
  PIN transducer_l15_csm_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 839.840 2500.000 840.440 ;
    END
  END transducer_l15_csm_data[28]
  PIN transducer_l15_csm_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END transducer_l15_csm_data[29]
  PIN transducer_l15_csm_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END transducer_l15_csm_data[2]
  PIN transducer_l15_csm_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.410 2496.000 1790.690 2500.000 ;
    END
  END transducer_l15_csm_data[30]
  PIN transducer_l15_csm_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 2496.000 261.190 2500.000 ;
    END
  END transducer_l15_csm_data[31]
  PIN transducer_l15_csm_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 2496.000 84.090 2500.000 ;
    END
  END transducer_l15_csm_data[32]
  PIN transducer_l15_csm_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 2496.000 644.370 2500.000 ;
    END
  END transducer_l15_csm_data[3]
  PIN transducer_l15_csm_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 2496.000 805.370 2500.000 ;
    END
  END transducer_l15_csm_data[4]
  PIN transducer_l15_csm_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 2496.000 844.010 2500.000 ;
    END
  END transducer_l15_csm_data[5]
  PIN transducer_l15_csm_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 0.000 1832.550 4.000 ;
    END
  END transducer_l15_csm_data[6]
  PIN transducer_l15_csm_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2332.440 4.000 2333.040 ;
    END
  END transducer_l15_csm_data[7]
  PIN transducer_l15_csm_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END transducer_l15_csm_data[8]
  PIN transducer_l15_csm_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END transducer_l15_csm_data[9]
  PIN transducer_l15_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 221.040 2500.000 221.640 ;
    END
  END transducer_l15_data[0]
  PIN transducer_l15_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 0.000 1835.770 4.000 ;
    END
  END transducer_l15_data[10]
  PIN transducer_l15_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END transducer_l15_data[11]
  PIN transducer_l15_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 2496.000 222.550 2500.000 ;
    END
  END transducer_l15_data[12]
  PIN transducer_l15_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1496.040 2500.000 1496.640 ;
    END
  END transducer_l15_data[13]
  PIN transducer_l15_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END transducer_l15_data[14]
  PIN transducer_l15_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END transducer_l15_data[15]
  PIN transducer_l15_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END transducer_l15_data[16]
  PIN transducer_l15_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 4.000 ;
    END
  END transducer_l15_data[17]
  PIN transducer_l15_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2424.240 4.000 2424.840 ;
    END
  END transducer_l15_data[18]
  PIN transducer_l15_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 258.440 2500.000 259.040 ;
    END
  END transducer_l15_data[19]
  PIN transducer_l15_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END transducer_l15_data[1]
  PIN transducer_l15_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 61.240 2500.000 61.840 ;
    END
  END transducer_l15_data[20]
  PIN transducer_l15_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 2496.000 2328.430 2500.000 ;
    END
  END transducer_l15_data[21]
  PIN transducer_l15_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 2496.000 1726.290 2500.000 ;
    END
  END transducer_l15_data[22]
  PIN transducer_l15_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 112.240 2500.000 112.840 ;
    END
  END transducer_l15_data[23]
  PIN transducer_l15_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END transducer_l15_data[24]
  PIN transducer_l15_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 860.240 2500.000 860.840 ;
    END
  END transducer_l15_data[25]
  PIN transducer_l15_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 2496.000 1909.830 2500.000 ;
    END
  END transducer_l15_data[26]
  PIN transducer_l15_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2135.240 4.000 2135.840 ;
    END
  END transducer_l15_data[27]
  PIN transducer_l15_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.030 2496.000 2341.310 2500.000 ;
    END
  END transducer_l15_data[28]
  PIN transducer_l15_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 27.240 2500.000 27.840 ;
    END
  END transducer_l15_data[29]
  PIN transducer_l15_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 2496.000 406.090 2500.000 ;
    END
  END transducer_l15_data[2]
  PIN transducer_l15_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1183.240 2500.000 1183.840 ;
    END
  END transducer_l15_data[30]
  PIN transducer_l15_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1965.240 4.000 1965.840 ;
    END
  END transducer_l15_data[31]
  PIN transducer_l15_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 564.440 2500.000 565.040 ;
    END
  END transducer_l15_data[32]
  PIN transducer_l15_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END transducer_l15_data[33]
  PIN transducer_l15_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END transducer_l15_data[34]
  PIN transducer_l15_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2495.640 2500.000 2496.240 ;
    END
  END transducer_l15_data[35]
  PIN transducer_l15_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 0.000 1829.330 4.000 ;
    END
  END transducer_l15_data[36]
  PIN transducer_l15_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.130 2496.000 2035.410 2500.000 ;
    END
  END transducer_l15_data[37]
  PIN transducer_l15_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END transducer_l15_data[38]
  PIN transducer_l15_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 581.440 2500.000 582.040 ;
    END
  END transducer_l15_data[39]
  PIN transducer_l15_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END transducer_l15_data[3]
  PIN transducer_l15_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 2496.000 560.650 2500.000 ;
    END
  END transducer_l15_data[40]
  PIN transducer_l15_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 2496.000 1768.150 2500.000 ;
    END
  END transducer_l15_data[41]
  PIN transducer_l15_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END transducer_l15_data[42]
  PIN transducer_l15_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END transducer_l15_data[43]
  PIN transducer_l15_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1271.640 2500.000 1272.240 ;
    END
  END transducer_l15_data[44]
  PIN transducer_l15_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END transducer_l15_data[45]
  PIN transducer_l15_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1815.640 2500.000 1816.240 ;
    END
  END transducer_l15_data[46]
  PIN transducer_l15_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 2496.000 93.750 2500.000 ;
    END
  END transducer_l15_data[47]
  PIN transducer_l15_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1931.240 4.000 1931.840 ;
    END
  END transducer_l15_data[48]
  PIN transducer_l15_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END transducer_l15_data[49]
  PIN transducer_l15_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END transducer_l15_data[4]
  PIN transducer_l15_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 0.000 1735.950 4.000 ;
    END
  END transducer_l15_data[50]
  PIN transducer_l15_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.910 2496.000 2032.190 2500.000 ;
    END
  END transducer_l15_data[51]
  PIN transducer_l15_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.330 2496.000 2228.610 2500.000 ;
    END
  END transducer_l15_data[52]
  PIN transducer_l15_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 0.000 1954.910 4.000 ;
    END
  END transducer_l15_data[53]
  PIN transducer_l15_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.050 2496.000 2473.330 2500.000 ;
    END
  END transducer_l15_data[54]
  PIN transducer_l15_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1587.840 2500.000 1588.440 ;
    END
  END transducer_l15_data[55]
  PIN transducer_l15_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 459.040 2500.000 459.640 ;
    END
  END transducer_l15_data[56]
  PIN transducer_l15_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END transducer_l15_data[57]
  PIN transducer_l15_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 2496.000 1124.150 2500.000 ;
    END
  END transducer_l15_data[58]
  PIN transducer_l15_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 4.000 ;
    END
  END transducer_l15_data[59]
  PIN transducer_l15_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.850 0.000 2441.130 4.000 ;
    END
  END transducer_l15_data[5]
  PIN transducer_l15_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1258.040 2500.000 1258.640 ;
    END
  END transducer_l15_data[60]
  PIN transducer_l15_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END transducer_l15_data[61]
  PIN transducer_l15_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 0.000 1632.910 4.000 ;
    END
  END transducer_l15_data[62]
  PIN transducer_l15_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END transducer_l15_data[63]
  PIN transducer_l15_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1968.640 4.000 1969.240 ;
    END
  END transducer_l15_data[6]
  PIN transducer_l15_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2301.840 2500.000 2302.440 ;
    END
  END transducer_l15_data[7]
  PIN transducer_l15_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 2496.000 1600.710 2500.000 ;
    END
  END transducer_l15_data[8]
  PIN transducer_l15_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END transducer_l15_data[9]
  PIN transducer_l15_data_next_entry[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 2496.000 901.970 2500.000 ;
    END
  END transducer_l15_data_next_entry[0]
  PIN transducer_l15_data_next_entry[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1757.840 2500.000 1758.440 ;
    END
  END transducer_l15_data_next_entry[10]
  PIN transducer_l15_data_next_entry[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.850 0.000 2280.130 4.000 ;
    END
  END transducer_l15_data_next_entry[11]
  PIN transducer_l15_data_next_entry[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 2496.000 885.870 2500.000 ;
    END
  END transducer_l15_data_next_entry[12]
  PIN transducer_l15_data_next_entry[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 0.000 2186.750 4.000 ;
    END
  END transducer_l15_data_next_entry[13]
  PIN transducer_l15_data_next_entry[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 4.000 ;
    END
  END transducer_l15_data_next_entry[14]
  PIN transducer_l15_data_next_entry[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END transducer_l15_data_next_entry[15]
  PIN transducer_l15_data_next_entry[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 408.040 2500.000 408.640 ;
    END
  END transducer_l15_data_next_entry[16]
  PIN transducer_l15_data_next_entry[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1220.640 2500.000 1221.240 ;
    END
  END transducer_l15_data_next_entry[17]
  PIN transducer_l15_data_next_entry[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2176.040 4.000 2176.640 ;
    END
  END transducer_l15_data_next_entry[18]
  PIN transducer_l15_data_next_entry[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 2496.000 2019.310 2500.000 ;
    END
  END transducer_l15_data_next_entry[19]
  PIN transducer_l15_data_next_entry[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END transducer_l15_data_next_entry[1]
  PIN transducer_l15_data_next_entry[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END transducer_l15_data_next_entry[20]
  PIN transducer_l15_data_next_entry[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END transducer_l15_data_next_entry[21]
  PIN transducer_l15_data_next_entry[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END transducer_l15_data_next_entry[22]
  PIN transducer_l15_data_next_entry[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END transducer_l15_data_next_entry[23]
  PIN transducer_l15_data_next_entry[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1887.040 2500.000 1887.640 ;
    END
  END transducer_l15_data_next_entry[24]
  PIN transducer_l15_data_next_entry[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 0.000 1623.250 4.000 ;
    END
  END transducer_l15_data_next_entry[25]
  PIN transducer_l15_data_next_entry[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 2496.000 889.090 2500.000 ;
    END
  END transducer_l15_data_next_entry[26]
  PIN transducer_l15_data_next_entry[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 2496.000 1581.390 2500.000 ;
    END
  END transducer_l15_data_next_entry[27]
  PIN transducer_l15_data_next_entry[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END transducer_l15_data_next_entry[28]
  PIN transducer_l15_data_next_entry[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END transducer_l15_data_next_entry[29]
  PIN transducer_l15_data_next_entry[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2060.440 2500.000 2061.040 ;
    END
  END transducer_l15_data_next_entry[2]
  PIN transducer_l15_data_next_entry[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 2496.000 1716.630 2500.000 ;
    END
  END transducer_l15_data_next_entry[30]
  PIN transducer_l15_data_next_entry[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END transducer_l15_data_next_entry[31]
  PIN transducer_l15_data_next_entry[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.170 2496.000 2460.450 2500.000 ;
    END
  END transducer_l15_data_next_entry[32]
  PIN transducer_l15_data_next_entry[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1217.240 2500.000 1217.840 ;
    END
  END transducer_l15_data_next_entry[33]
  PIN transducer_l15_data_next_entry[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.330 0.000 1906.610 4.000 ;
    END
  END transducer_l15_data_next_entry[34]
  PIN transducer_l15_data_next_entry[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 2496.000 1455.810 2500.000 ;
    END
  END transducer_l15_data_next_entry[35]
  PIN transducer_l15_data_next_entry[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2352.840 4.000 2353.440 ;
    END
  END transducer_l15_data_next_entry[36]
  PIN transducer_l15_data_next_entry[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END transducer_l15_data_next_entry[37]
  PIN transducer_l15_data_next_entry[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1968.640 2500.000 1969.240 ;
    END
  END transducer_l15_data_next_entry[38]
  PIN transducer_l15_data_next_entry[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.330 0.000 2228.610 4.000 ;
    END
  END transducer_l15_data_next_entry[39]
  PIN transducer_l15_data_next_entry[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1064.240 2500.000 1064.840 ;
    END
  END transducer_l15_data_next_entry[3]
  PIN transducer_l15_data_next_entry[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END transducer_l15_data_next_entry[40]
  PIN transducer_l15_data_next_entry[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 312.840 2500.000 313.440 ;
    END
  END transducer_l15_data_next_entry[41]
  PIN transducer_l15_data_next_entry[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END transducer_l15_data_next_entry[42]
  PIN transducer_l15_data_next_entry[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 0.000 1336.670 4.000 ;
    END
  END transducer_l15_data_next_entry[43]
  PIN transducer_l15_data_next_entry[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1407.640 2500.000 1408.240 ;
    END
  END transducer_l15_data_next_entry[44]
  PIN transducer_l15_data_next_entry[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 2496.000 1497.670 2500.000 ;
    END
  END transducer_l15_data_next_entry[45]
  PIN transducer_l15_data_next_entry[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.370 2496.000 2331.650 2500.000 ;
    END
  END transducer_l15_data_next_entry[46]
  PIN transducer_l15_data_next_entry[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 309.440 2500.000 310.040 ;
    END
  END transducer_l15_data_next_entry[47]
  PIN transducer_l15_data_next_entry[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END transducer_l15_data_next_entry[48]
  PIN transducer_l15_data_next_entry[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1740.840 2500.000 1741.440 ;
    END
  END transducer_l15_data_next_entry[49]
  PIN transducer_l15_data_next_entry[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END transducer_l15_data_next_entry[4]
  PIN transducer_l15_data_next_entry[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.710 2496.000 2321.990 2500.000 ;
    END
  END transducer_l15_data_next_entry[50]
  PIN transducer_l15_data_next_entry[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 2496.000 1484.790 2500.000 ;
    END
  END transducer_l15_data_next_entry[51]
  PIN transducer_l15_data_next_entry[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 452.240 2500.000 452.840 ;
    END
  END transducer_l15_data_next_entry[52]
  PIN transducer_l15_data_next_entry[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 2496.000 1420.390 2500.000 ;
    END
  END transducer_l15_data_next_entry[53]
  PIN transducer_l15_data_next_entry[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 0.000 1764.930 4.000 ;
    END
  END transducer_l15_data_next_entry[54]
  PIN transducer_l15_data_next_entry[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END transducer_l15_data_next_entry[55]
  PIN transducer_l15_data_next_entry[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.770 0.000 1752.050 4.000 ;
    END
  END transducer_l15_data_next_entry[56]
  PIN transducer_l15_data_next_entry[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END transducer_l15_data_next_entry[57]
  PIN transducer_l15_data_next_entry[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.790 0.000 2045.070 4.000 ;
    END
  END transducer_l15_data_next_entry[58]
  PIN transducer_l15_data_next_entry[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END transducer_l15_data_next_entry[59]
  PIN transducer_l15_data_next_entry[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1798.640 4.000 1799.240 ;
    END
  END transducer_l15_data_next_entry[5]
  PIN transducer_l15_data_next_entry[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 2496.000 396.430 2500.000 ;
    END
  END transducer_l15_data_next_entry[60]
  PIN transducer_l15_data_next_entry[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END transducer_l15_data_next_entry[61]
  PIN transducer_l15_data_next_entry[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END transducer_l15_data_next_entry[62]
  PIN transducer_l15_data_next_entry[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END transducer_l15_data_next_entry[63]
  PIN transducer_l15_data_next_entry[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 2496.000 1075.850 2500.000 ;
    END
  END transducer_l15_data_next_entry[6]
  PIN transducer_l15_data_next_entry[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 2496.000 518.790 2500.000 ;
    END
  END transducer_l15_data_next_entry[7]
  PIN transducer_l15_data_next_entry[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 0.000 1378.530 4.000 ;
    END
  END transducer_l15_data_next_entry[8]
  PIN transducer_l15_data_next_entry[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 2496.000 1549.190 2500.000 ;
    END
  END transducer_l15_data_next_entry[9]
  PIN transducer_l15_invalidate_cacheline
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 771.840 2500.000 772.440 ;
    END
  END transducer_l15_invalidate_cacheline
  PIN transducer_l15_l1rplway[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END transducer_l15_l1rplway[0]
  PIN transducer_l15_l1rplway[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2057.040 2500.000 2057.640 ;
    END
  END transducer_l15_l1rplway[1]
  PIN transducer_l15_nc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END transducer_l15_nc
  PIN transducer_l15_prefetch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END transducer_l15_prefetch
  PIN transducer_l15_req_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END transducer_l15_req_ack
  PIN transducer_l15_rqtype[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1927.840 2500.000 1928.440 ;
    END
  END transducer_l15_rqtype[0]
  PIN transducer_l15_rqtype[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 0.000 1513.770 4.000 ;
    END
  END transducer_l15_rqtype[1]
  PIN transducer_l15_rqtype[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 2496.000 1571.730 2500.000 ;
    END
  END transducer_l15_rqtype[2]
  PIN transducer_l15_rqtype[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 2496.000 1552.410 2500.000 ;
    END
  END transducer_l15_rqtype[3]
  PIN transducer_l15_rqtype[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2281.440 4.000 2282.040 ;
    END
  END transducer_l15_rqtype[4]
  PIN transducer_l15_size[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 2496.000 251.530 2500.000 ;
    END
  END transducer_l15_size[0]
  PIN transducer_l15_size[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.750 0.000 1781.030 4.000 ;
    END
  END transducer_l15_size[1]
  PIN transducer_l15_size[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END transducer_l15_size[2]
  PIN transducer_l15_threadid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2094.440 4.000 2095.040 ;
    END
  END transducer_l15_threadid
  PIN transducer_l15_val
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1210.440 2500.000 1211.040 ;
    END
  END transducer_l15_val
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 2489.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 2494.360 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 2494.360 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 2494.360 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 2494.360 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 2494.360 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 792.630 2494.360 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 945.810 2494.360 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1098.990 2494.360 1100.590 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1252.170 2494.360 1253.770 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1405.350 2494.360 1406.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1558.530 2494.360 1560.130 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1711.710 2494.360 1713.310 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1864.890 2494.360 1866.490 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2018.070 2494.360 2019.670 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2171.250 2494.360 2172.850 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2324.430 2494.360 2326.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2477.610 2494.360 2479.210 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2489.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 2489.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 103.320 2494.360 104.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 256.500 2494.360 258.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 409.680 2494.360 411.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 562.860 2494.360 564.460 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 716.040 2494.360 717.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 869.220 2494.360 870.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1022.400 2494.360 1024.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1175.580 2494.360 1177.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1328.760 2494.360 1330.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1481.940 2494.360 1483.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1635.120 2494.360 1636.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1788.300 2494.360 1789.900 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1941.480 2494.360 1943.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2094.660 2494.360 2096.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2247.840 2494.360 2249.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2401.020 2494.360 2402.620 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2494.120 2488.885 ;
      LAYER met1 ;
        RECT 0.070 5.820 2499.110 2490.120 ;
      LAYER met2 ;
        RECT 0.650 2495.720 3.030 2499.525 ;
        RECT 3.870 2495.720 6.250 2499.525 ;
        RECT 7.090 2495.720 9.470 2499.525 ;
        RECT 10.310 2495.720 12.690 2499.525 ;
        RECT 13.530 2495.720 15.910 2499.525 ;
        RECT 16.750 2495.720 19.130 2499.525 ;
        RECT 19.970 2495.720 22.350 2499.525 ;
        RECT 23.190 2495.720 25.570 2499.525 ;
        RECT 26.410 2495.720 28.790 2499.525 ;
        RECT 29.630 2495.720 32.010 2499.525 ;
        RECT 32.850 2495.720 35.230 2499.525 ;
        RECT 36.070 2495.720 41.670 2499.525 ;
        RECT 42.510 2495.720 44.890 2499.525 ;
        RECT 45.730 2495.720 48.110 2499.525 ;
        RECT 48.950 2495.720 51.330 2499.525 ;
        RECT 52.170 2495.720 54.550 2499.525 ;
        RECT 55.390 2495.720 57.770 2499.525 ;
        RECT 58.610 2495.720 60.990 2499.525 ;
        RECT 61.830 2495.720 64.210 2499.525 ;
        RECT 65.050 2495.720 67.430 2499.525 ;
        RECT 68.270 2495.720 70.650 2499.525 ;
        RECT 71.490 2495.720 73.870 2499.525 ;
        RECT 74.710 2495.720 77.090 2499.525 ;
        RECT 77.930 2495.720 80.310 2499.525 ;
        RECT 81.150 2495.720 83.530 2499.525 ;
        RECT 84.370 2495.720 86.750 2499.525 ;
        RECT 87.590 2495.720 93.190 2499.525 ;
        RECT 94.030 2495.720 96.410 2499.525 ;
        RECT 97.250 2495.720 99.630 2499.525 ;
        RECT 100.470 2495.720 102.850 2499.525 ;
        RECT 103.690 2495.720 106.070 2499.525 ;
        RECT 106.910 2495.720 109.290 2499.525 ;
        RECT 110.130 2495.720 112.510 2499.525 ;
        RECT 113.350 2495.720 115.730 2499.525 ;
        RECT 116.570 2495.720 118.950 2499.525 ;
        RECT 119.790 2495.720 122.170 2499.525 ;
        RECT 123.010 2495.720 125.390 2499.525 ;
        RECT 126.230 2495.720 128.610 2499.525 ;
        RECT 129.450 2495.720 131.830 2499.525 ;
        RECT 132.670 2495.720 135.050 2499.525 ;
        RECT 135.890 2495.720 138.270 2499.525 ;
        RECT 139.110 2495.720 144.710 2499.525 ;
        RECT 145.550 2495.720 147.930 2499.525 ;
        RECT 148.770 2495.720 151.150 2499.525 ;
        RECT 151.990 2495.720 154.370 2499.525 ;
        RECT 155.210 2495.720 157.590 2499.525 ;
        RECT 158.430 2495.720 160.810 2499.525 ;
        RECT 161.650 2495.720 164.030 2499.525 ;
        RECT 164.870 2495.720 167.250 2499.525 ;
        RECT 168.090 2495.720 170.470 2499.525 ;
        RECT 171.310 2495.720 173.690 2499.525 ;
        RECT 174.530 2495.720 176.910 2499.525 ;
        RECT 177.750 2495.720 180.130 2499.525 ;
        RECT 180.970 2495.720 183.350 2499.525 ;
        RECT 184.190 2495.720 186.570 2499.525 ;
        RECT 187.410 2495.720 189.790 2499.525 ;
        RECT 190.630 2495.720 196.230 2499.525 ;
        RECT 197.070 2495.720 199.450 2499.525 ;
        RECT 200.290 2495.720 202.670 2499.525 ;
        RECT 203.510 2495.720 205.890 2499.525 ;
        RECT 206.730 2495.720 209.110 2499.525 ;
        RECT 209.950 2495.720 212.330 2499.525 ;
        RECT 213.170 2495.720 215.550 2499.525 ;
        RECT 216.390 2495.720 218.770 2499.525 ;
        RECT 219.610 2495.720 221.990 2499.525 ;
        RECT 222.830 2495.720 225.210 2499.525 ;
        RECT 226.050 2495.720 228.430 2499.525 ;
        RECT 229.270 2495.720 231.650 2499.525 ;
        RECT 232.490 2495.720 234.870 2499.525 ;
        RECT 235.710 2495.720 238.090 2499.525 ;
        RECT 238.930 2495.720 241.310 2499.525 ;
        RECT 242.150 2495.720 247.750 2499.525 ;
        RECT 248.590 2495.720 250.970 2499.525 ;
        RECT 251.810 2495.720 254.190 2499.525 ;
        RECT 255.030 2495.720 257.410 2499.525 ;
        RECT 258.250 2495.720 260.630 2499.525 ;
        RECT 261.470 2495.720 263.850 2499.525 ;
        RECT 264.690 2495.720 267.070 2499.525 ;
        RECT 267.910 2495.720 270.290 2499.525 ;
        RECT 271.130 2495.720 273.510 2499.525 ;
        RECT 274.350 2495.720 276.730 2499.525 ;
        RECT 277.570 2495.720 279.950 2499.525 ;
        RECT 280.790 2495.720 283.170 2499.525 ;
        RECT 284.010 2495.720 286.390 2499.525 ;
        RECT 287.230 2495.720 289.610 2499.525 ;
        RECT 290.450 2495.720 292.830 2499.525 ;
        RECT 293.670 2495.720 299.270 2499.525 ;
        RECT 300.110 2495.720 302.490 2499.525 ;
        RECT 303.330 2495.720 305.710 2499.525 ;
        RECT 306.550 2495.720 308.930 2499.525 ;
        RECT 309.770 2495.720 312.150 2499.525 ;
        RECT 312.990 2495.720 315.370 2499.525 ;
        RECT 316.210 2495.720 318.590 2499.525 ;
        RECT 319.430 2495.720 321.810 2499.525 ;
        RECT 322.650 2495.720 325.030 2499.525 ;
        RECT 325.870 2495.720 328.250 2499.525 ;
        RECT 329.090 2495.720 331.470 2499.525 ;
        RECT 332.310 2495.720 334.690 2499.525 ;
        RECT 335.530 2495.720 337.910 2499.525 ;
        RECT 338.750 2495.720 341.130 2499.525 ;
        RECT 341.970 2495.720 344.350 2499.525 ;
        RECT 345.190 2495.720 350.790 2499.525 ;
        RECT 351.630 2495.720 354.010 2499.525 ;
        RECT 354.850 2495.720 357.230 2499.525 ;
        RECT 358.070 2495.720 360.450 2499.525 ;
        RECT 361.290 2495.720 363.670 2499.525 ;
        RECT 364.510 2495.720 366.890 2499.525 ;
        RECT 367.730 2495.720 370.110 2499.525 ;
        RECT 370.950 2495.720 373.330 2499.525 ;
        RECT 374.170 2495.720 376.550 2499.525 ;
        RECT 377.390 2495.720 379.770 2499.525 ;
        RECT 380.610 2495.720 382.990 2499.525 ;
        RECT 383.830 2495.720 386.210 2499.525 ;
        RECT 387.050 2495.720 389.430 2499.525 ;
        RECT 390.270 2495.720 392.650 2499.525 ;
        RECT 393.490 2495.720 395.870 2499.525 ;
        RECT 396.710 2495.720 402.310 2499.525 ;
        RECT 403.150 2495.720 405.530 2499.525 ;
        RECT 406.370 2495.720 408.750 2499.525 ;
        RECT 409.590 2495.720 411.970 2499.525 ;
        RECT 412.810 2495.720 415.190 2499.525 ;
        RECT 416.030 2495.720 418.410 2499.525 ;
        RECT 419.250 2495.720 421.630 2499.525 ;
        RECT 422.470 2495.720 424.850 2499.525 ;
        RECT 425.690 2495.720 428.070 2499.525 ;
        RECT 428.910 2495.720 431.290 2499.525 ;
        RECT 432.130 2495.720 434.510 2499.525 ;
        RECT 435.350 2495.720 437.730 2499.525 ;
        RECT 438.570 2495.720 440.950 2499.525 ;
        RECT 441.790 2495.720 444.170 2499.525 ;
        RECT 445.010 2495.720 450.610 2499.525 ;
        RECT 451.450 2495.720 453.830 2499.525 ;
        RECT 454.670 2495.720 457.050 2499.525 ;
        RECT 457.890 2495.720 460.270 2499.525 ;
        RECT 461.110 2495.720 463.490 2499.525 ;
        RECT 464.330 2495.720 466.710 2499.525 ;
        RECT 467.550 2495.720 469.930 2499.525 ;
        RECT 470.770 2495.720 473.150 2499.525 ;
        RECT 473.990 2495.720 476.370 2499.525 ;
        RECT 477.210 2495.720 479.590 2499.525 ;
        RECT 480.430 2495.720 482.810 2499.525 ;
        RECT 483.650 2495.720 486.030 2499.525 ;
        RECT 486.870 2495.720 489.250 2499.525 ;
        RECT 490.090 2495.720 492.470 2499.525 ;
        RECT 493.310 2495.720 495.690 2499.525 ;
        RECT 496.530 2495.720 502.130 2499.525 ;
        RECT 502.970 2495.720 505.350 2499.525 ;
        RECT 506.190 2495.720 508.570 2499.525 ;
        RECT 509.410 2495.720 511.790 2499.525 ;
        RECT 512.630 2495.720 515.010 2499.525 ;
        RECT 515.850 2495.720 518.230 2499.525 ;
        RECT 519.070 2495.720 521.450 2499.525 ;
        RECT 522.290 2495.720 524.670 2499.525 ;
        RECT 525.510 2495.720 527.890 2499.525 ;
        RECT 528.730 2495.720 531.110 2499.525 ;
        RECT 531.950 2495.720 534.330 2499.525 ;
        RECT 535.170 2495.720 537.550 2499.525 ;
        RECT 538.390 2495.720 540.770 2499.525 ;
        RECT 541.610 2495.720 543.990 2499.525 ;
        RECT 544.830 2495.720 547.210 2499.525 ;
        RECT 548.050 2495.720 553.650 2499.525 ;
        RECT 554.490 2495.720 556.870 2499.525 ;
        RECT 557.710 2495.720 560.090 2499.525 ;
        RECT 560.930 2495.720 563.310 2499.525 ;
        RECT 564.150 2495.720 566.530 2499.525 ;
        RECT 567.370 2495.720 569.750 2499.525 ;
        RECT 570.590 2495.720 572.970 2499.525 ;
        RECT 573.810 2495.720 576.190 2499.525 ;
        RECT 577.030 2495.720 579.410 2499.525 ;
        RECT 580.250 2495.720 582.630 2499.525 ;
        RECT 583.470 2495.720 585.850 2499.525 ;
        RECT 586.690 2495.720 589.070 2499.525 ;
        RECT 589.910 2495.720 592.290 2499.525 ;
        RECT 593.130 2495.720 595.510 2499.525 ;
        RECT 596.350 2495.720 598.730 2499.525 ;
        RECT 599.570 2495.720 605.170 2499.525 ;
        RECT 606.010 2495.720 608.390 2499.525 ;
        RECT 609.230 2495.720 611.610 2499.525 ;
        RECT 612.450 2495.720 614.830 2499.525 ;
        RECT 615.670 2495.720 618.050 2499.525 ;
        RECT 618.890 2495.720 621.270 2499.525 ;
        RECT 622.110 2495.720 624.490 2499.525 ;
        RECT 625.330 2495.720 627.710 2499.525 ;
        RECT 628.550 2495.720 630.930 2499.525 ;
        RECT 631.770 2495.720 634.150 2499.525 ;
        RECT 634.990 2495.720 637.370 2499.525 ;
        RECT 638.210 2495.720 640.590 2499.525 ;
        RECT 641.430 2495.720 643.810 2499.525 ;
        RECT 644.650 2495.720 647.030 2499.525 ;
        RECT 647.870 2495.720 650.250 2499.525 ;
        RECT 651.090 2495.720 656.690 2499.525 ;
        RECT 657.530 2495.720 659.910 2499.525 ;
        RECT 660.750 2495.720 663.130 2499.525 ;
        RECT 663.970 2495.720 666.350 2499.525 ;
        RECT 667.190 2495.720 669.570 2499.525 ;
        RECT 670.410 2495.720 672.790 2499.525 ;
        RECT 673.630 2495.720 676.010 2499.525 ;
        RECT 676.850 2495.720 679.230 2499.525 ;
        RECT 680.070 2495.720 682.450 2499.525 ;
        RECT 683.290 2495.720 685.670 2499.525 ;
        RECT 686.510 2495.720 688.890 2499.525 ;
        RECT 689.730 2495.720 692.110 2499.525 ;
        RECT 692.950 2495.720 695.330 2499.525 ;
        RECT 696.170 2495.720 698.550 2499.525 ;
        RECT 699.390 2495.720 701.770 2499.525 ;
        RECT 702.610 2495.720 708.210 2499.525 ;
        RECT 709.050 2495.720 711.430 2499.525 ;
        RECT 712.270 2495.720 714.650 2499.525 ;
        RECT 715.490 2495.720 717.870 2499.525 ;
        RECT 718.710 2495.720 721.090 2499.525 ;
        RECT 721.930 2495.720 724.310 2499.525 ;
        RECT 725.150 2495.720 727.530 2499.525 ;
        RECT 728.370 2495.720 730.750 2499.525 ;
        RECT 731.590 2495.720 733.970 2499.525 ;
        RECT 734.810 2495.720 737.190 2499.525 ;
        RECT 738.030 2495.720 740.410 2499.525 ;
        RECT 741.250 2495.720 743.630 2499.525 ;
        RECT 744.470 2495.720 746.850 2499.525 ;
        RECT 747.690 2495.720 750.070 2499.525 ;
        RECT 750.910 2495.720 753.290 2499.525 ;
        RECT 754.130 2495.720 759.730 2499.525 ;
        RECT 760.570 2495.720 762.950 2499.525 ;
        RECT 763.790 2495.720 766.170 2499.525 ;
        RECT 767.010 2495.720 769.390 2499.525 ;
        RECT 770.230 2495.720 772.610 2499.525 ;
        RECT 773.450 2495.720 775.830 2499.525 ;
        RECT 776.670 2495.720 779.050 2499.525 ;
        RECT 779.890 2495.720 782.270 2499.525 ;
        RECT 783.110 2495.720 785.490 2499.525 ;
        RECT 786.330 2495.720 788.710 2499.525 ;
        RECT 789.550 2495.720 791.930 2499.525 ;
        RECT 792.770 2495.720 795.150 2499.525 ;
        RECT 795.990 2495.720 798.370 2499.525 ;
        RECT 799.210 2495.720 801.590 2499.525 ;
        RECT 802.430 2495.720 804.810 2499.525 ;
        RECT 805.650 2495.720 811.250 2499.525 ;
        RECT 812.090 2495.720 814.470 2499.525 ;
        RECT 815.310 2495.720 817.690 2499.525 ;
        RECT 818.530 2495.720 820.910 2499.525 ;
        RECT 821.750 2495.720 824.130 2499.525 ;
        RECT 824.970 2495.720 827.350 2499.525 ;
        RECT 828.190 2495.720 830.570 2499.525 ;
        RECT 831.410 2495.720 833.790 2499.525 ;
        RECT 834.630 2495.720 837.010 2499.525 ;
        RECT 837.850 2495.720 840.230 2499.525 ;
        RECT 841.070 2495.720 843.450 2499.525 ;
        RECT 844.290 2495.720 846.670 2499.525 ;
        RECT 847.510 2495.720 849.890 2499.525 ;
        RECT 850.730 2495.720 853.110 2499.525 ;
        RECT 853.950 2495.720 856.330 2499.525 ;
        RECT 857.170 2495.720 862.770 2499.525 ;
        RECT 863.610 2495.720 865.990 2499.525 ;
        RECT 866.830 2495.720 869.210 2499.525 ;
        RECT 870.050 2495.720 872.430 2499.525 ;
        RECT 873.270 2495.720 875.650 2499.525 ;
        RECT 876.490 2495.720 878.870 2499.525 ;
        RECT 879.710 2495.720 882.090 2499.525 ;
        RECT 882.930 2495.720 885.310 2499.525 ;
        RECT 886.150 2495.720 888.530 2499.525 ;
        RECT 889.370 2495.720 891.750 2499.525 ;
        RECT 892.590 2495.720 894.970 2499.525 ;
        RECT 895.810 2495.720 898.190 2499.525 ;
        RECT 899.030 2495.720 901.410 2499.525 ;
        RECT 902.250 2495.720 904.630 2499.525 ;
        RECT 905.470 2495.720 907.850 2499.525 ;
        RECT 908.690 2495.720 914.290 2499.525 ;
        RECT 915.130 2495.720 917.510 2499.525 ;
        RECT 918.350 2495.720 920.730 2499.525 ;
        RECT 921.570 2495.720 923.950 2499.525 ;
        RECT 924.790 2495.720 927.170 2499.525 ;
        RECT 928.010 2495.720 930.390 2499.525 ;
        RECT 931.230 2495.720 933.610 2499.525 ;
        RECT 934.450 2495.720 936.830 2499.525 ;
        RECT 937.670 2495.720 940.050 2499.525 ;
        RECT 940.890 2495.720 943.270 2499.525 ;
        RECT 944.110 2495.720 946.490 2499.525 ;
        RECT 947.330 2495.720 949.710 2499.525 ;
        RECT 950.550 2495.720 952.930 2499.525 ;
        RECT 953.770 2495.720 956.150 2499.525 ;
        RECT 956.990 2495.720 959.370 2499.525 ;
        RECT 960.210 2495.720 965.810 2499.525 ;
        RECT 966.650 2495.720 969.030 2499.525 ;
        RECT 969.870 2495.720 972.250 2499.525 ;
        RECT 973.090 2495.720 975.470 2499.525 ;
        RECT 976.310 2495.720 978.690 2499.525 ;
        RECT 979.530 2495.720 981.910 2499.525 ;
        RECT 982.750 2495.720 985.130 2499.525 ;
        RECT 985.970 2495.720 988.350 2499.525 ;
        RECT 989.190 2495.720 991.570 2499.525 ;
        RECT 992.410 2495.720 994.790 2499.525 ;
        RECT 995.630 2495.720 998.010 2499.525 ;
        RECT 998.850 2495.720 1001.230 2499.525 ;
        RECT 1002.070 2495.720 1004.450 2499.525 ;
        RECT 1005.290 2495.720 1007.670 2499.525 ;
        RECT 1008.510 2495.720 1010.890 2499.525 ;
        RECT 1011.730 2495.720 1017.330 2499.525 ;
        RECT 1018.170 2495.720 1020.550 2499.525 ;
        RECT 1021.390 2495.720 1023.770 2499.525 ;
        RECT 1024.610 2495.720 1026.990 2499.525 ;
        RECT 1027.830 2495.720 1030.210 2499.525 ;
        RECT 1031.050 2495.720 1033.430 2499.525 ;
        RECT 1034.270 2495.720 1036.650 2499.525 ;
        RECT 1037.490 2495.720 1039.870 2499.525 ;
        RECT 1040.710 2495.720 1043.090 2499.525 ;
        RECT 1043.930 2495.720 1046.310 2499.525 ;
        RECT 1047.150 2495.720 1049.530 2499.525 ;
        RECT 1050.370 2495.720 1052.750 2499.525 ;
        RECT 1053.590 2495.720 1055.970 2499.525 ;
        RECT 1056.810 2495.720 1059.190 2499.525 ;
        RECT 1060.030 2495.720 1062.410 2499.525 ;
        RECT 1063.250 2495.720 1068.850 2499.525 ;
        RECT 1069.690 2495.720 1072.070 2499.525 ;
        RECT 1072.910 2495.720 1075.290 2499.525 ;
        RECT 1076.130 2495.720 1078.510 2499.525 ;
        RECT 1079.350 2495.720 1081.730 2499.525 ;
        RECT 1082.570 2495.720 1084.950 2499.525 ;
        RECT 1085.790 2495.720 1088.170 2499.525 ;
        RECT 1089.010 2495.720 1091.390 2499.525 ;
        RECT 1092.230 2495.720 1094.610 2499.525 ;
        RECT 1095.450 2495.720 1097.830 2499.525 ;
        RECT 1098.670 2495.720 1101.050 2499.525 ;
        RECT 1101.890 2495.720 1104.270 2499.525 ;
        RECT 1105.110 2495.720 1107.490 2499.525 ;
        RECT 1108.330 2495.720 1110.710 2499.525 ;
        RECT 1111.550 2495.720 1117.150 2499.525 ;
        RECT 1117.990 2495.720 1120.370 2499.525 ;
        RECT 1121.210 2495.720 1123.590 2499.525 ;
        RECT 1124.430 2495.720 1126.810 2499.525 ;
        RECT 1127.650 2495.720 1130.030 2499.525 ;
        RECT 1130.870 2495.720 1133.250 2499.525 ;
        RECT 1134.090 2495.720 1136.470 2499.525 ;
        RECT 1137.310 2495.720 1139.690 2499.525 ;
        RECT 1140.530 2495.720 1142.910 2499.525 ;
        RECT 1143.750 2495.720 1146.130 2499.525 ;
        RECT 1146.970 2495.720 1149.350 2499.525 ;
        RECT 1150.190 2495.720 1152.570 2499.525 ;
        RECT 1153.410 2495.720 1155.790 2499.525 ;
        RECT 1156.630 2495.720 1159.010 2499.525 ;
        RECT 1159.850 2495.720 1162.230 2499.525 ;
        RECT 1163.070 2495.720 1168.670 2499.525 ;
        RECT 1169.510 2495.720 1171.890 2499.525 ;
        RECT 1172.730 2495.720 1175.110 2499.525 ;
        RECT 1175.950 2495.720 1178.330 2499.525 ;
        RECT 1179.170 2495.720 1181.550 2499.525 ;
        RECT 1182.390 2495.720 1184.770 2499.525 ;
        RECT 1185.610 2495.720 1187.990 2499.525 ;
        RECT 1188.830 2495.720 1191.210 2499.525 ;
        RECT 1192.050 2495.720 1194.430 2499.525 ;
        RECT 1195.270 2495.720 1197.650 2499.525 ;
        RECT 1198.490 2495.720 1200.870 2499.525 ;
        RECT 1201.710 2495.720 1204.090 2499.525 ;
        RECT 1204.930 2495.720 1207.310 2499.525 ;
        RECT 1208.150 2495.720 1210.530 2499.525 ;
        RECT 1211.370 2495.720 1213.750 2499.525 ;
        RECT 1214.590 2495.720 1220.190 2499.525 ;
        RECT 1221.030 2495.720 1223.410 2499.525 ;
        RECT 1224.250 2495.720 1226.630 2499.525 ;
        RECT 1227.470 2495.720 1229.850 2499.525 ;
        RECT 1230.690 2495.720 1233.070 2499.525 ;
        RECT 1233.910 2495.720 1236.290 2499.525 ;
        RECT 1237.130 2495.720 1239.510 2499.525 ;
        RECT 1240.350 2495.720 1242.730 2499.525 ;
        RECT 1243.570 2495.720 1245.950 2499.525 ;
        RECT 1246.790 2495.720 1249.170 2499.525 ;
        RECT 1250.010 2495.720 1252.390 2499.525 ;
        RECT 1253.230 2495.720 1255.610 2499.525 ;
        RECT 1256.450 2495.720 1258.830 2499.525 ;
        RECT 1259.670 2495.720 1262.050 2499.525 ;
        RECT 1262.890 2495.720 1265.270 2499.525 ;
        RECT 1266.110 2495.720 1271.710 2499.525 ;
        RECT 1272.550 2495.720 1274.930 2499.525 ;
        RECT 1275.770 2495.720 1278.150 2499.525 ;
        RECT 1278.990 2495.720 1281.370 2499.525 ;
        RECT 1282.210 2495.720 1284.590 2499.525 ;
        RECT 1285.430 2495.720 1287.810 2499.525 ;
        RECT 1288.650 2495.720 1291.030 2499.525 ;
        RECT 1291.870 2495.720 1294.250 2499.525 ;
        RECT 1295.090 2495.720 1297.470 2499.525 ;
        RECT 1298.310 2495.720 1300.690 2499.525 ;
        RECT 1301.530 2495.720 1303.910 2499.525 ;
        RECT 1304.750 2495.720 1307.130 2499.525 ;
        RECT 1307.970 2495.720 1310.350 2499.525 ;
        RECT 1311.190 2495.720 1313.570 2499.525 ;
        RECT 1314.410 2495.720 1316.790 2499.525 ;
        RECT 1317.630 2495.720 1323.230 2499.525 ;
        RECT 1324.070 2495.720 1326.450 2499.525 ;
        RECT 1327.290 2495.720 1329.670 2499.525 ;
        RECT 1330.510 2495.720 1332.890 2499.525 ;
        RECT 1333.730 2495.720 1336.110 2499.525 ;
        RECT 1336.950 2495.720 1339.330 2499.525 ;
        RECT 1340.170 2495.720 1342.550 2499.525 ;
        RECT 1343.390 2495.720 1345.770 2499.525 ;
        RECT 1346.610 2495.720 1348.990 2499.525 ;
        RECT 1349.830 2495.720 1352.210 2499.525 ;
        RECT 1353.050 2495.720 1355.430 2499.525 ;
        RECT 1356.270 2495.720 1358.650 2499.525 ;
        RECT 1359.490 2495.720 1361.870 2499.525 ;
        RECT 1362.710 2495.720 1365.090 2499.525 ;
        RECT 1365.930 2495.720 1368.310 2499.525 ;
        RECT 1369.150 2495.720 1374.750 2499.525 ;
        RECT 1375.590 2495.720 1377.970 2499.525 ;
        RECT 1378.810 2495.720 1381.190 2499.525 ;
        RECT 1382.030 2495.720 1384.410 2499.525 ;
        RECT 1385.250 2495.720 1387.630 2499.525 ;
        RECT 1388.470 2495.720 1390.850 2499.525 ;
        RECT 1391.690 2495.720 1394.070 2499.525 ;
        RECT 1394.910 2495.720 1397.290 2499.525 ;
        RECT 1398.130 2495.720 1400.510 2499.525 ;
        RECT 1401.350 2495.720 1403.730 2499.525 ;
        RECT 1404.570 2495.720 1406.950 2499.525 ;
        RECT 1407.790 2495.720 1410.170 2499.525 ;
        RECT 1411.010 2495.720 1413.390 2499.525 ;
        RECT 1414.230 2495.720 1416.610 2499.525 ;
        RECT 1417.450 2495.720 1419.830 2499.525 ;
        RECT 1420.670 2495.720 1426.270 2499.525 ;
        RECT 1427.110 2495.720 1429.490 2499.525 ;
        RECT 1430.330 2495.720 1432.710 2499.525 ;
        RECT 1433.550 2495.720 1435.930 2499.525 ;
        RECT 1436.770 2495.720 1439.150 2499.525 ;
        RECT 1439.990 2495.720 1442.370 2499.525 ;
        RECT 1443.210 2495.720 1445.590 2499.525 ;
        RECT 1446.430 2495.720 1448.810 2499.525 ;
        RECT 1449.650 2495.720 1452.030 2499.525 ;
        RECT 1452.870 2495.720 1455.250 2499.525 ;
        RECT 1456.090 2495.720 1458.470 2499.525 ;
        RECT 1459.310 2495.720 1461.690 2499.525 ;
        RECT 1462.530 2495.720 1464.910 2499.525 ;
        RECT 1465.750 2495.720 1468.130 2499.525 ;
        RECT 1468.970 2495.720 1471.350 2499.525 ;
        RECT 1472.190 2495.720 1477.790 2499.525 ;
        RECT 1478.630 2495.720 1481.010 2499.525 ;
        RECT 1481.850 2495.720 1484.230 2499.525 ;
        RECT 1485.070 2495.720 1487.450 2499.525 ;
        RECT 1488.290 2495.720 1490.670 2499.525 ;
        RECT 1491.510 2495.720 1493.890 2499.525 ;
        RECT 1494.730 2495.720 1497.110 2499.525 ;
        RECT 1497.950 2495.720 1500.330 2499.525 ;
        RECT 1501.170 2495.720 1503.550 2499.525 ;
        RECT 1504.390 2495.720 1506.770 2499.525 ;
        RECT 1507.610 2495.720 1509.990 2499.525 ;
        RECT 1510.830 2495.720 1513.210 2499.525 ;
        RECT 1514.050 2495.720 1516.430 2499.525 ;
        RECT 1517.270 2495.720 1519.650 2499.525 ;
        RECT 1520.490 2495.720 1522.870 2499.525 ;
        RECT 1523.710 2495.720 1529.310 2499.525 ;
        RECT 1530.150 2495.720 1532.530 2499.525 ;
        RECT 1533.370 2495.720 1535.750 2499.525 ;
        RECT 1536.590 2495.720 1538.970 2499.525 ;
        RECT 1539.810 2495.720 1542.190 2499.525 ;
        RECT 1543.030 2495.720 1545.410 2499.525 ;
        RECT 1546.250 2495.720 1548.630 2499.525 ;
        RECT 1549.470 2495.720 1551.850 2499.525 ;
        RECT 1552.690 2495.720 1555.070 2499.525 ;
        RECT 1555.910 2495.720 1558.290 2499.525 ;
        RECT 1559.130 2495.720 1561.510 2499.525 ;
        RECT 1562.350 2495.720 1564.730 2499.525 ;
        RECT 1565.570 2495.720 1567.950 2499.525 ;
        RECT 1568.790 2495.720 1571.170 2499.525 ;
        RECT 1572.010 2495.720 1574.390 2499.525 ;
        RECT 1575.230 2495.720 1580.830 2499.525 ;
        RECT 1581.670 2495.720 1584.050 2499.525 ;
        RECT 1584.890 2495.720 1587.270 2499.525 ;
        RECT 1588.110 2495.720 1590.490 2499.525 ;
        RECT 1591.330 2495.720 1593.710 2499.525 ;
        RECT 1594.550 2495.720 1596.930 2499.525 ;
        RECT 1597.770 2495.720 1600.150 2499.525 ;
        RECT 1600.990 2495.720 1603.370 2499.525 ;
        RECT 1604.210 2495.720 1606.590 2499.525 ;
        RECT 1607.430 2495.720 1609.810 2499.525 ;
        RECT 1610.650 2495.720 1613.030 2499.525 ;
        RECT 1613.870 2495.720 1616.250 2499.525 ;
        RECT 1617.090 2495.720 1619.470 2499.525 ;
        RECT 1620.310 2495.720 1622.690 2499.525 ;
        RECT 1623.530 2495.720 1625.910 2499.525 ;
        RECT 1626.750 2495.720 1632.350 2499.525 ;
        RECT 1633.190 2495.720 1635.570 2499.525 ;
        RECT 1636.410 2495.720 1638.790 2499.525 ;
        RECT 1639.630 2495.720 1642.010 2499.525 ;
        RECT 1642.850 2495.720 1645.230 2499.525 ;
        RECT 1646.070 2495.720 1648.450 2499.525 ;
        RECT 1649.290 2495.720 1651.670 2499.525 ;
        RECT 1652.510 2495.720 1654.890 2499.525 ;
        RECT 1655.730 2495.720 1658.110 2499.525 ;
        RECT 1658.950 2495.720 1661.330 2499.525 ;
        RECT 1662.170 2495.720 1664.550 2499.525 ;
        RECT 1665.390 2495.720 1667.770 2499.525 ;
        RECT 1668.610 2495.720 1670.990 2499.525 ;
        RECT 1671.830 2495.720 1674.210 2499.525 ;
        RECT 1675.050 2495.720 1677.430 2499.525 ;
        RECT 1678.270 2495.720 1683.870 2499.525 ;
        RECT 1684.710 2495.720 1687.090 2499.525 ;
        RECT 1687.930 2495.720 1690.310 2499.525 ;
        RECT 1691.150 2495.720 1693.530 2499.525 ;
        RECT 1694.370 2495.720 1696.750 2499.525 ;
        RECT 1697.590 2495.720 1699.970 2499.525 ;
        RECT 1700.810 2495.720 1703.190 2499.525 ;
        RECT 1704.030 2495.720 1706.410 2499.525 ;
        RECT 1707.250 2495.720 1709.630 2499.525 ;
        RECT 1710.470 2495.720 1712.850 2499.525 ;
        RECT 1713.690 2495.720 1716.070 2499.525 ;
        RECT 1716.910 2495.720 1719.290 2499.525 ;
        RECT 1720.130 2495.720 1722.510 2499.525 ;
        RECT 1723.350 2495.720 1725.730 2499.525 ;
        RECT 1726.570 2495.720 1728.950 2499.525 ;
        RECT 1729.790 2495.720 1735.390 2499.525 ;
        RECT 1736.230 2495.720 1738.610 2499.525 ;
        RECT 1739.450 2495.720 1741.830 2499.525 ;
        RECT 1742.670 2495.720 1745.050 2499.525 ;
        RECT 1745.890 2495.720 1748.270 2499.525 ;
        RECT 1749.110 2495.720 1751.490 2499.525 ;
        RECT 1752.330 2495.720 1754.710 2499.525 ;
        RECT 1755.550 2495.720 1757.930 2499.525 ;
        RECT 1758.770 2495.720 1761.150 2499.525 ;
        RECT 1761.990 2495.720 1764.370 2499.525 ;
        RECT 1765.210 2495.720 1767.590 2499.525 ;
        RECT 1768.430 2495.720 1770.810 2499.525 ;
        RECT 1771.650 2495.720 1774.030 2499.525 ;
        RECT 1774.870 2495.720 1777.250 2499.525 ;
        RECT 1778.090 2495.720 1780.470 2499.525 ;
        RECT 1781.310 2495.720 1786.910 2499.525 ;
        RECT 1787.750 2495.720 1790.130 2499.525 ;
        RECT 1790.970 2495.720 1793.350 2499.525 ;
        RECT 1794.190 2495.720 1796.570 2499.525 ;
        RECT 1797.410 2495.720 1799.790 2499.525 ;
        RECT 1800.630 2495.720 1803.010 2499.525 ;
        RECT 1803.850 2495.720 1806.230 2499.525 ;
        RECT 1807.070 2495.720 1809.450 2499.525 ;
        RECT 1810.290 2495.720 1812.670 2499.525 ;
        RECT 1813.510 2495.720 1815.890 2499.525 ;
        RECT 1816.730 2495.720 1819.110 2499.525 ;
        RECT 1819.950 2495.720 1822.330 2499.525 ;
        RECT 1823.170 2495.720 1825.550 2499.525 ;
        RECT 1826.390 2495.720 1828.770 2499.525 ;
        RECT 1829.610 2495.720 1835.210 2499.525 ;
        RECT 1836.050 2495.720 1838.430 2499.525 ;
        RECT 1839.270 2495.720 1841.650 2499.525 ;
        RECT 1842.490 2495.720 1844.870 2499.525 ;
        RECT 1845.710 2495.720 1848.090 2499.525 ;
        RECT 1848.930 2495.720 1851.310 2499.525 ;
        RECT 1852.150 2495.720 1854.530 2499.525 ;
        RECT 1855.370 2495.720 1857.750 2499.525 ;
        RECT 1858.590 2495.720 1860.970 2499.525 ;
        RECT 1861.810 2495.720 1864.190 2499.525 ;
        RECT 1865.030 2495.720 1867.410 2499.525 ;
        RECT 1868.250 2495.720 1870.630 2499.525 ;
        RECT 1871.470 2495.720 1873.850 2499.525 ;
        RECT 1874.690 2495.720 1877.070 2499.525 ;
        RECT 1877.910 2495.720 1880.290 2499.525 ;
        RECT 1881.130 2495.720 1886.730 2499.525 ;
        RECT 1887.570 2495.720 1889.950 2499.525 ;
        RECT 1890.790 2495.720 1893.170 2499.525 ;
        RECT 1894.010 2495.720 1896.390 2499.525 ;
        RECT 1897.230 2495.720 1899.610 2499.525 ;
        RECT 1900.450 2495.720 1902.830 2499.525 ;
        RECT 1903.670 2495.720 1906.050 2499.525 ;
        RECT 1906.890 2495.720 1909.270 2499.525 ;
        RECT 1910.110 2495.720 1912.490 2499.525 ;
        RECT 1913.330 2495.720 1915.710 2499.525 ;
        RECT 1916.550 2495.720 1918.930 2499.525 ;
        RECT 1919.770 2495.720 1922.150 2499.525 ;
        RECT 1922.990 2495.720 1925.370 2499.525 ;
        RECT 1926.210 2495.720 1928.590 2499.525 ;
        RECT 1929.430 2495.720 1931.810 2499.525 ;
        RECT 1932.650 2495.720 1938.250 2499.525 ;
        RECT 1939.090 2495.720 1941.470 2499.525 ;
        RECT 1942.310 2495.720 1944.690 2499.525 ;
        RECT 1945.530 2495.720 1947.910 2499.525 ;
        RECT 1948.750 2495.720 1951.130 2499.525 ;
        RECT 1951.970 2495.720 1954.350 2499.525 ;
        RECT 1955.190 2495.720 1957.570 2499.525 ;
        RECT 1958.410 2495.720 1960.790 2499.525 ;
        RECT 1961.630 2495.720 1964.010 2499.525 ;
        RECT 1964.850 2495.720 1967.230 2499.525 ;
        RECT 1968.070 2495.720 1970.450 2499.525 ;
        RECT 1971.290 2495.720 1973.670 2499.525 ;
        RECT 1974.510 2495.720 1976.890 2499.525 ;
        RECT 1977.730 2495.720 1980.110 2499.525 ;
        RECT 1980.950 2495.720 1983.330 2499.525 ;
        RECT 1984.170 2495.720 1989.770 2499.525 ;
        RECT 1990.610 2495.720 1992.990 2499.525 ;
        RECT 1993.830 2495.720 1996.210 2499.525 ;
        RECT 1997.050 2495.720 1999.430 2499.525 ;
        RECT 2000.270 2495.720 2002.650 2499.525 ;
        RECT 2003.490 2495.720 2005.870 2499.525 ;
        RECT 2006.710 2495.720 2009.090 2499.525 ;
        RECT 2009.930 2495.720 2012.310 2499.525 ;
        RECT 2013.150 2495.720 2015.530 2499.525 ;
        RECT 2016.370 2495.720 2018.750 2499.525 ;
        RECT 2019.590 2495.720 2021.970 2499.525 ;
        RECT 2022.810 2495.720 2025.190 2499.525 ;
        RECT 2026.030 2495.720 2028.410 2499.525 ;
        RECT 2029.250 2495.720 2031.630 2499.525 ;
        RECT 2032.470 2495.720 2034.850 2499.525 ;
        RECT 2035.690 2495.720 2041.290 2499.525 ;
        RECT 2042.130 2495.720 2044.510 2499.525 ;
        RECT 2045.350 2495.720 2047.730 2499.525 ;
        RECT 2048.570 2495.720 2050.950 2499.525 ;
        RECT 2051.790 2495.720 2054.170 2499.525 ;
        RECT 2055.010 2495.720 2057.390 2499.525 ;
        RECT 2058.230 2495.720 2060.610 2499.525 ;
        RECT 2061.450 2495.720 2063.830 2499.525 ;
        RECT 2064.670 2495.720 2067.050 2499.525 ;
        RECT 2067.890 2495.720 2070.270 2499.525 ;
        RECT 2071.110 2495.720 2073.490 2499.525 ;
        RECT 2074.330 2495.720 2076.710 2499.525 ;
        RECT 2077.550 2495.720 2079.930 2499.525 ;
        RECT 2080.770 2495.720 2083.150 2499.525 ;
        RECT 2083.990 2495.720 2086.370 2499.525 ;
        RECT 2087.210 2495.720 2092.810 2499.525 ;
        RECT 2093.650 2495.720 2096.030 2499.525 ;
        RECT 2096.870 2495.720 2099.250 2499.525 ;
        RECT 2100.090 2495.720 2102.470 2499.525 ;
        RECT 2103.310 2495.720 2105.690 2499.525 ;
        RECT 2106.530 2495.720 2108.910 2499.525 ;
        RECT 2109.750 2495.720 2112.130 2499.525 ;
        RECT 2112.970 2495.720 2115.350 2499.525 ;
        RECT 2116.190 2495.720 2118.570 2499.525 ;
        RECT 2119.410 2495.720 2121.790 2499.525 ;
        RECT 2122.630 2495.720 2125.010 2499.525 ;
        RECT 2125.850 2495.720 2128.230 2499.525 ;
        RECT 2129.070 2495.720 2131.450 2499.525 ;
        RECT 2132.290 2495.720 2134.670 2499.525 ;
        RECT 2135.510 2495.720 2137.890 2499.525 ;
        RECT 2138.730 2495.720 2144.330 2499.525 ;
        RECT 2145.170 2495.720 2147.550 2499.525 ;
        RECT 2148.390 2495.720 2150.770 2499.525 ;
        RECT 2151.610 2495.720 2153.990 2499.525 ;
        RECT 2154.830 2495.720 2157.210 2499.525 ;
        RECT 2158.050 2495.720 2160.430 2499.525 ;
        RECT 2161.270 2495.720 2163.650 2499.525 ;
        RECT 2164.490 2495.720 2166.870 2499.525 ;
        RECT 2167.710 2495.720 2170.090 2499.525 ;
        RECT 2170.930 2495.720 2173.310 2499.525 ;
        RECT 2174.150 2495.720 2176.530 2499.525 ;
        RECT 2177.370 2495.720 2179.750 2499.525 ;
        RECT 2180.590 2495.720 2182.970 2499.525 ;
        RECT 2183.810 2495.720 2186.190 2499.525 ;
        RECT 2187.030 2495.720 2189.410 2499.525 ;
        RECT 2190.250 2495.720 2195.850 2499.525 ;
        RECT 2196.690 2495.720 2199.070 2499.525 ;
        RECT 2199.910 2495.720 2202.290 2499.525 ;
        RECT 2203.130 2495.720 2205.510 2499.525 ;
        RECT 2206.350 2495.720 2208.730 2499.525 ;
        RECT 2209.570 2495.720 2211.950 2499.525 ;
        RECT 2212.790 2495.720 2215.170 2499.525 ;
        RECT 2216.010 2495.720 2218.390 2499.525 ;
        RECT 2219.230 2495.720 2221.610 2499.525 ;
        RECT 2222.450 2495.720 2224.830 2499.525 ;
        RECT 2225.670 2495.720 2228.050 2499.525 ;
        RECT 2228.890 2495.720 2231.270 2499.525 ;
        RECT 2232.110 2495.720 2234.490 2499.525 ;
        RECT 2235.330 2495.720 2237.710 2499.525 ;
        RECT 2238.550 2495.720 2240.930 2499.525 ;
        RECT 2241.770 2495.720 2247.370 2499.525 ;
        RECT 2248.210 2495.720 2250.590 2499.525 ;
        RECT 2251.430 2495.720 2253.810 2499.525 ;
        RECT 2254.650 2495.720 2257.030 2499.525 ;
        RECT 2257.870 2495.720 2260.250 2499.525 ;
        RECT 2261.090 2495.720 2263.470 2499.525 ;
        RECT 2264.310 2495.720 2266.690 2499.525 ;
        RECT 2267.530 2495.720 2269.910 2499.525 ;
        RECT 2270.750 2495.720 2273.130 2499.525 ;
        RECT 2273.970 2495.720 2276.350 2499.525 ;
        RECT 2277.190 2495.720 2279.570 2499.525 ;
        RECT 2280.410 2495.720 2282.790 2499.525 ;
        RECT 2283.630 2495.720 2286.010 2499.525 ;
        RECT 2286.850 2495.720 2289.230 2499.525 ;
        RECT 2290.070 2495.720 2292.450 2499.525 ;
        RECT 2293.290 2495.720 2298.890 2499.525 ;
        RECT 2299.730 2495.720 2302.110 2499.525 ;
        RECT 2302.950 2495.720 2305.330 2499.525 ;
        RECT 2306.170 2495.720 2308.550 2499.525 ;
        RECT 2309.390 2495.720 2311.770 2499.525 ;
        RECT 2312.610 2495.720 2314.990 2499.525 ;
        RECT 2315.830 2495.720 2318.210 2499.525 ;
        RECT 2319.050 2495.720 2321.430 2499.525 ;
        RECT 2322.270 2495.720 2324.650 2499.525 ;
        RECT 2325.490 2495.720 2327.870 2499.525 ;
        RECT 2328.710 2495.720 2331.090 2499.525 ;
        RECT 2331.930 2495.720 2334.310 2499.525 ;
        RECT 2335.150 2495.720 2337.530 2499.525 ;
        RECT 2338.370 2495.720 2340.750 2499.525 ;
        RECT 2341.590 2495.720 2343.970 2499.525 ;
        RECT 2344.810 2495.720 2350.410 2499.525 ;
        RECT 2351.250 2495.720 2353.630 2499.525 ;
        RECT 2354.470 2495.720 2356.850 2499.525 ;
        RECT 2357.690 2495.720 2360.070 2499.525 ;
        RECT 2360.910 2495.720 2363.290 2499.525 ;
        RECT 2364.130 2495.720 2366.510 2499.525 ;
        RECT 2367.350 2495.720 2369.730 2499.525 ;
        RECT 2370.570 2495.720 2372.950 2499.525 ;
        RECT 2373.790 2495.720 2376.170 2499.525 ;
        RECT 2377.010 2495.720 2379.390 2499.525 ;
        RECT 2380.230 2495.720 2382.610 2499.525 ;
        RECT 2383.450 2495.720 2385.830 2499.525 ;
        RECT 2386.670 2495.720 2389.050 2499.525 ;
        RECT 2389.890 2495.720 2392.270 2499.525 ;
        RECT 2393.110 2495.720 2395.490 2499.525 ;
        RECT 2396.330 2495.720 2401.930 2499.525 ;
        RECT 2402.770 2495.720 2405.150 2499.525 ;
        RECT 2405.990 2495.720 2408.370 2499.525 ;
        RECT 2409.210 2495.720 2411.590 2499.525 ;
        RECT 2412.430 2495.720 2414.810 2499.525 ;
        RECT 2415.650 2495.720 2418.030 2499.525 ;
        RECT 2418.870 2495.720 2421.250 2499.525 ;
        RECT 2422.090 2495.720 2424.470 2499.525 ;
        RECT 2425.310 2495.720 2427.690 2499.525 ;
        RECT 2428.530 2495.720 2430.910 2499.525 ;
        RECT 2431.750 2495.720 2434.130 2499.525 ;
        RECT 2434.970 2495.720 2437.350 2499.525 ;
        RECT 2438.190 2495.720 2440.570 2499.525 ;
        RECT 2441.410 2495.720 2443.790 2499.525 ;
        RECT 2444.630 2495.720 2447.010 2499.525 ;
        RECT 2447.850 2495.720 2453.450 2499.525 ;
        RECT 2454.290 2495.720 2456.670 2499.525 ;
        RECT 2457.510 2495.720 2459.890 2499.525 ;
        RECT 2460.730 2495.720 2463.110 2499.525 ;
        RECT 2463.950 2495.720 2466.330 2499.525 ;
        RECT 2467.170 2495.720 2469.550 2499.525 ;
        RECT 2470.390 2495.720 2472.770 2499.525 ;
        RECT 2473.610 2495.720 2475.990 2499.525 ;
        RECT 2476.830 2495.720 2479.210 2499.525 ;
        RECT 2480.050 2495.720 2482.430 2499.525 ;
        RECT 2483.270 2495.720 2485.650 2499.525 ;
        RECT 2486.490 2495.720 2488.870 2499.525 ;
        RECT 2489.710 2495.720 2492.090 2499.525 ;
        RECT 2492.930 2495.720 2495.310 2499.525 ;
        RECT 2496.150 2495.720 2498.530 2499.525 ;
        RECT 0.100 4.280 2499.080 2495.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
        RECT 148.770 0.155 154.370 4.280 ;
        RECT 155.210 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 167.250 4.280 ;
        RECT 168.090 0.155 170.470 4.280 ;
        RECT 171.310 0.155 173.690 4.280 ;
        RECT 174.530 0.155 176.910 4.280 ;
        RECT 177.750 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 186.570 4.280 ;
        RECT 187.410 0.155 189.790 4.280 ;
        RECT 190.630 0.155 193.010 4.280 ;
        RECT 193.850 0.155 196.230 4.280 ;
        RECT 197.070 0.155 199.450 4.280 ;
        RECT 200.290 0.155 205.890 4.280 ;
        RECT 206.730 0.155 209.110 4.280 ;
        RECT 209.950 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.550 4.280 ;
        RECT 216.390 0.155 218.770 4.280 ;
        RECT 219.610 0.155 221.990 4.280 ;
        RECT 222.830 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 231.650 4.280 ;
        RECT 232.490 0.155 234.870 4.280 ;
        RECT 235.710 0.155 238.090 4.280 ;
        RECT 238.930 0.155 241.310 4.280 ;
        RECT 242.150 0.155 244.530 4.280 ;
        RECT 245.370 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 257.410 4.280 ;
        RECT 258.250 0.155 260.630 4.280 ;
        RECT 261.470 0.155 263.850 4.280 ;
        RECT 264.690 0.155 267.070 4.280 ;
        RECT 267.910 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 276.730 4.280 ;
        RECT 277.570 0.155 279.950 4.280 ;
        RECT 280.790 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 308.930 4.280 ;
        RECT 309.770 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 334.690 4.280 ;
        RECT 335.530 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 350.790 4.280 ;
        RECT 351.630 0.155 354.010 4.280 ;
        RECT 354.850 0.155 360.450 4.280 ;
        RECT 361.290 0.155 363.670 4.280 ;
        RECT 364.510 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 373.330 4.280 ;
        RECT 374.170 0.155 376.550 4.280 ;
        RECT 377.390 0.155 379.770 4.280 ;
        RECT 380.610 0.155 382.990 4.280 ;
        RECT 383.830 0.155 386.210 4.280 ;
        RECT 387.050 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 395.870 4.280 ;
        RECT 396.710 0.155 399.090 4.280 ;
        RECT 399.930 0.155 402.310 4.280 ;
        RECT 403.150 0.155 405.530 4.280 ;
        RECT 406.370 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 418.410 4.280 ;
        RECT 419.250 0.155 421.630 4.280 ;
        RECT 422.470 0.155 424.850 4.280 ;
        RECT 425.690 0.155 428.070 4.280 ;
        RECT 428.910 0.155 431.290 4.280 ;
        RECT 432.130 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 440.950 4.280 ;
        RECT 441.790 0.155 444.170 4.280 ;
        RECT 445.010 0.155 447.390 4.280 ;
        RECT 448.230 0.155 450.610 4.280 ;
        RECT 451.450 0.155 453.830 4.280 ;
        RECT 454.670 0.155 457.050 4.280 ;
        RECT 457.890 0.155 463.490 4.280 ;
        RECT 464.330 0.155 466.710 4.280 ;
        RECT 467.550 0.155 469.930 4.280 ;
        RECT 470.770 0.155 473.150 4.280 ;
        RECT 473.990 0.155 476.370 4.280 ;
        RECT 477.210 0.155 479.590 4.280 ;
        RECT 480.430 0.155 482.810 4.280 ;
        RECT 483.650 0.155 486.030 4.280 ;
        RECT 486.870 0.155 489.250 4.280 ;
        RECT 490.090 0.155 492.470 4.280 ;
        RECT 493.310 0.155 495.690 4.280 ;
        RECT 496.530 0.155 498.910 4.280 ;
        RECT 499.750 0.155 502.130 4.280 ;
        RECT 502.970 0.155 505.350 4.280 ;
        RECT 506.190 0.155 508.570 4.280 ;
        RECT 509.410 0.155 515.010 4.280 ;
        RECT 515.850 0.155 518.230 4.280 ;
        RECT 519.070 0.155 521.450 4.280 ;
        RECT 522.290 0.155 524.670 4.280 ;
        RECT 525.510 0.155 527.890 4.280 ;
        RECT 528.730 0.155 531.110 4.280 ;
        RECT 531.950 0.155 534.330 4.280 ;
        RECT 535.170 0.155 537.550 4.280 ;
        RECT 538.390 0.155 540.770 4.280 ;
        RECT 541.610 0.155 543.990 4.280 ;
        RECT 544.830 0.155 547.210 4.280 ;
        RECT 548.050 0.155 550.430 4.280 ;
        RECT 551.270 0.155 553.650 4.280 ;
        RECT 554.490 0.155 556.870 4.280 ;
        RECT 557.710 0.155 560.090 4.280 ;
        RECT 560.930 0.155 566.530 4.280 ;
        RECT 567.370 0.155 569.750 4.280 ;
        RECT 570.590 0.155 572.970 4.280 ;
        RECT 573.810 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 582.630 4.280 ;
        RECT 583.470 0.155 585.850 4.280 ;
        RECT 586.690 0.155 589.070 4.280 ;
        RECT 589.910 0.155 592.290 4.280 ;
        RECT 593.130 0.155 595.510 4.280 ;
        RECT 596.350 0.155 598.730 4.280 ;
        RECT 599.570 0.155 601.950 4.280 ;
        RECT 602.790 0.155 605.170 4.280 ;
        RECT 606.010 0.155 608.390 4.280 ;
        RECT 609.230 0.155 611.610 4.280 ;
        RECT 612.450 0.155 618.050 4.280 ;
        RECT 618.890 0.155 621.270 4.280 ;
        RECT 622.110 0.155 624.490 4.280 ;
        RECT 625.330 0.155 627.710 4.280 ;
        RECT 628.550 0.155 630.930 4.280 ;
        RECT 631.770 0.155 634.150 4.280 ;
        RECT 634.990 0.155 637.370 4.280 ;
        RECT 638.210 0.155 640.590 4.280 ;
        RECT 641.430 0.155 643.810 4.280 ;
        RECT 644.650 0.155 647.030 4.280 ;
        RECT 647.870 0.155 650.250 4.280 ;
        RECT 651.090 0.155 653.470 4.280 ;
        RECT 654.310 0.155 656.690 4.280 ;
        RECT 657.530 0.155 659.910 4.280 ;
        RECT 660.750 0.155 663.130 4.280 ;
        RECT 663.970 0.155 669.570 4.280 ;
        RECT 670.410 0.155 672.790 4.280 ;
        RECT 673.630 0.155 676.010 4.280 ;
        RECT 676.850 0.155 679.230 4.280 ;
        RECT 680.070 0.155 682.450 4.280 ;
        RECT 683.290 0.155 685.670 4.280 ;
        RECT 686.510 0.155 688.890 4.280 ;
        RECT 689.730 0.155 692.110 4.280 ;
        RECT 692.950 0.155 695.330 4.280 ;
        RECT 696.170 0.155 698.550 4.280 ;
        RECT 699.390 0.155 701.770 4.280 ;
        RECT 702.610 0.155 704.990 4.280 ;
        RECT 705.830 0.155 708.210 4.280 ;
        RECT 709.050 0.155 711.430 4.280 ;
        RECT 712.270 0.155 717.870 4.280 ;
        RECT 718.710 0.155 721.090 4.280 ;
        RECT 721.930 0.155 724.310 4.280 ;
        RECT 725.150 0.155 727.530 4.280 ;
        RECT 728.370 0.155 730.750 4.280 ;
        RECT 731.590 0.155 733.970 4.280 ;
        RECT 734.810 0.155 737.190 4.280 ;
        RECT 738.030 0.155 740.410 4.280 ;
        RECT 741.250 0.155 743.630 4.280 ;
        RECT 744.470 0.155 746.850 4.280 ;
        RECT 747.690 0.155 750.070 4.280 ;
        RECT 750.910 0.155 753.290 4.280 ;
        RECT 754.130 0.155 756.510 4.280 ;
        RECT 757.350 0.155 759.730 4.280 ;
        RECT 760.570 0.155 762.950 4.280 ;
        RECT 763.790 0.155 769.390 4.280 ;
        RECT 770.230 0.155 772.610 4.280 ;
        RECT 773.450 0.155 775.830 4.280 ;
        RECT 776.670 0.155 779.050 4.280 ;
        RECT 779.890 0.155 782.270 4.280 ;
        RECT 783.110 0.155 785.490 4.280 ;
        RECT 786.330 0.155 788.710 4.280 ;
        RECT 789.550 0.155 791.930 4.280 ;
        RECT 792.770 0.155 795.150 4.280 ;
        RECT 795.990 0.155 798.370 4.280 ;
        RECT 799.210 0.155 801.590 4.280 ;
        RECT 802.430 0.155 804.810 4.280 ;
        RECT 805.650 0.155 808.030 4.280 ;
        RECT 808.870 0.155 811.250 4.280 ;
        RECT 812.090 0.155 814.470 4.280 ;
        RECT 815.310 0.155 820.910 4.280 ;
        RECT 821.750 0.155 824.130 4.280 ;
        RECT 824.970 0.155 827.350 4.280 ;
        RECT 828.190 0.155 830.570 4.280 ;
        RECT 831.410 0.155 833.790 4.280 ;
        RECT 834.630 0.155 837.010 4.280 ;
        RECT 837.850 0.155 840.230 4.280 ;
        RECT 841.070 0.155 843.450 4.280 ;
        RECT 844.290 0.155 846.670 4.280 ;
        RECT 847.510 0.155 849.890 4.280 ;
        RECT 850.730 0.155 853.110 4.280 ;
        RECT 853.950 0.155 856.330 4.280 ;
        RECT 857.170 0.155 859.550 4.280 ;
        RECT 860.390 0.155 862.770 4.280 ;
        RECT 863.610 0.155 865.990 4.280 ;
        RECT 866.830 0.155 872.430 4.280 ;
        RECT 873.270 0.155 875.650 4.280 ;
        RECT 876.490 0.155 878.870 4.280 ;
        RECT 879.710 0.155 882.090 4.280 ;
        RECT 882.930 0.155 885.310 4.280 ;
        RECT 886.150 0.155 888.530 4.280 ;
        RECT 889.370 0.155 891.750 4.280 ;
        RECT 892.590 0.155 894.970 4.280 ;
        RECT 895.810 0.155 898.190 4.280 ;
        RECT 899.030 0.155 901.410 4.280 ;
        RECT 902.250 0.155 904.630 4.280 ;
        RECT 905.470 0.155 907.850 4.280 ;
        RECT 908.690 0.155 911.070 4.280 ;
        RECT 911.910 0.155 914.290 4.280 ;
        RECT 915.130 0.155 917.510 4.280 ;
        RECT 918.350 0.155 923.950 4.280 ;
        RECT 924.790 0.155 927.170 4.280 ;
        RECT 928.010 0.155 930.390 4.280 ;
        RECT 931.230 0.155 933.610 4.280 ;
        RECT 934.450 0.155 936.830 4.280 ;
        RECT 937.670 0.155 940.050 4.280 ;
        RECT 940.890 0.155 943.270 4.280 ;
        RECT 944.110 0.155 946.490 4.280 ;
        RECT 947.330 0.155 949.710 4.280 ;
        RECT 950.550 0.155 952.930 4.280 ;
        RECT 953.770 0.155 956.150 4.280 ;
        RECT 956.990 0.155 959.370 4.280 ;
        RECT 960.210 0.155 962.590 4.280 ;
        RECT 963.430 0.155 965.810 4.280 ;
        RECT 966.650 0.155 969.030 4.280 ;
        RECT 969.870 0.155 975.470 4.280 ;
        RECT 976.310 0.155 978.690 4.280 ;
        RECT 979.530 0.155 981.910 4.280 ;
        RECT 982.750 0.155 985.130 4.280 ;
        RECT 985.970 0.155 988.350 4.280 ;
        RECT 989.190 0.155 991.570 4.280 ;
        RECT 992.410 0.155 994.790 4.280 ;
        RECT 995.630 0.155 998.010 4.280 ;
        RECT 998.850 0.155 1001.230 4.280 ;
        RECT 1002.070 0.155 1004.450 4.280 ;
        RECT 1005.290 0.155 1007.670 4.280 ;
        RECT 1008.510 0.155 1010.890 4.280 ;
        RECT 1011.730 0.155 1014.110 4.280 ;
        RECT 1014.950 0.155 1017.330 4.280 ;
        RECT 1018.170 0.155 1020.550 4.280 ;
        RECT 1021.390 0.155 1026.990 4.280 ;
        RECT 1027.830 0.155 1030.210 4.280 ;
        RECT 1031.050 0.155 1033.430 4.280 ;
        RECT 1034.270 0.155 1036.650 4.280 ;
        RECT 1037.490 0.155 1039.870 4.280 ;
        RECT 1040.710 0.155 1043.090 4.280 ;
        RECT 1043.930 0.155 1046.310 4.280 ;
        RECT 1047.150 0.155 1049.530 4.280 ;
        RECT 1050.370 0.155 1052.750 4.280 ;
        RECT 1053.590 0.155 1055.970 4.280 ;
        RECT 1056.810 0.155 1059.190 4.280 ;
        RECT 1060.030 0.155 1062.410 4.280 ;
        RECT 1063.250 0.155 1065.630 4.280 ;
        RECT 1066.470 0.155 1068.850 4.280 ;
        RECT 1069.690 0.155 1072.070 4.280 ;
        RECT 1072.910 0.155 1078.510 4.280 ;
        RECT 1079.350 0.155 1081.730 4.280 ;
        RECT 1082.570 0.155 1084.950 4.280 ;
        RECT 1085.790 0.155 1088.170 4.280 ;
        RECT 1089.010 0.155 1091.390 4.280 ;
        RECT 1092.230 0.155 1094.610 4.280 ;
        RECT 1095.450 0.155 1097.830 4.280 ;
        RECT 1098.670 0.155 1101.050 4.280 ;
        RECT 1101.890 0.155 1104.270 4.280 ;
        RECT 1105.110 0.155 1107.490 4.280 ;
        RECT 1108.330 0.155 1110.710 4.280 ;
        RECT 1111.550 0.155 1113.930 4.280 ;
        RECT 1114.770 0.155 1117.150 4.280 ;
        RECT 1117.990 0.155 1120.370 4.280 ;
        RECT 1121.210 0.155 1123.590 4.280 ;
        RECT 1124.430 0.155 1130.030 4.280 ;
        RECT 1130.870 0.155 1133.250 4.280 ;
        RECT 1134.090 0.155 1136.470 4.280 ;
        RECT 1137.310 0.155 1139.690 4.280 ;
        RECT 1140.530 0.155 1142.910 4.280 ;
        RECT 1143.750 0.155 1146.130 4.280 ;
        RECT 1146.970 0.155 1149.350 4.280 ;
        RECT 1150.190 0.155 1152.570 4.280 ;
        RECT 1153.410 0.155 1155.790 4.280 ;
        RECT 1156.630 0.155 1159.010 4.280 ;
        RECT 1159.850 0.155 1162.230 4.280 ;
        RECT 1163.070 0.155 1165.450 4.280 ;
        RECT 1166.290 0.155 1168.670 4.280 ;
        RECT 1169.510 0.155 1171.890 4.280 ;
        RECT 1172.730 0.155 1175.110 4.280 ;
        RECT 1175.950 0.155 1181.550 4.280 ;
        RECT 1182.390 0.155 1184.770 4.280 ;
        RECT 1185.610 0.155 1187.990 4.280 ;
        RECT 1188.830 0.155 1191.210 4.280 ;
        RECT 1192.050 0.155 1194.430 4.280 ;
        RECT 1195.270 0.155 1197.650 4.280 ;
        RECT 1198.490 0.155 1200.870 4.280 ;
        RECT 1201.710 0.155 1204.090 4.280 ;
        RECT 1204.930 0.155 1207.310 4.280 ;
        RECT 1208.150 0.155 1210.530 4.280 ;
        RECT 1211.370 0.155 1213.750 4.280 ;
        RECT 1214.590 0.155 1216.970 4.280 ;
        RECT 1217.810 0.155 1220.190 4.280 ;
        RECT 1221.030 0.155 1223.410 4.280 ;
        RECT 1224.250 0.155 1226.630 4.280 ;
        RECT 1227.470 0.155 1233.070 4.280 ;
        RECT 1233.910 0.155 1236.290 4.280 ;
        RECT 1237.130 0.155 1239.510 4.280 ;
        RECT 1240.350 0.155 1242.730 4.280 ;
        RECT 1243.570 0.155 1245.950 4.280 ;
        RECT 1246.790 0.155 1249.170 4.280 ;
        RECT 1250.010 0.155 1252.390 4.280 ;
        RECT 1253.230 0.155 1255.610 4.280 ;
        RECT 1256.450 0.155 1258.830 4.280 ;
        RECT 1259.670 0.155 1262.050 4.280 ;
        RECT 1262.890 0.155 1265.270 4.280 ;
        RECT 1266.110 0.155 1268.490 4.280 ;
        RECT 1269.330 0.155 1271.710 4.280 ;
        RECT 1272.550 0.155 1274.930 4.280 ;
        RECT 1275.770 0.155 1278.150 4.280 ;
        RECT 1278.990 0.155 1284.590 4.280 ;
        RECT 1285.430 0.155 1287.810 4.280 ;
        RECT 1288.650 0.155 1291.030 4.280 ;
        RECT 1291.870 0.155 1294.250 4.280 ;
        RECT 1295.090 0.155 1297.470 4.280 ;
        RECT 1298.310 0.155 1300.690 4.280 ;
        RECT 1301.530 0.155 1303.910 4.280 ;
        RECT 1304.750 0.155 1307.130 4.280 ;
        RECT 1307.970 0.155 1310.350 4.280 ;
        RECT 1311.190 0.155 1313.570 4.280 ;
        RECT 1314.410 0.155 1316.790 4.280 ;
        RECT 1317.630 0.155 1320.010 4.280 ;
        RECT 1320.850 0.155 1323.230 4.280 ;
        RECT 1324.070 0.155 1326.450 4.280 ;
        RECT 1327.290 0.155 1329.670 4.280 ;
        RECT 1330.510 0.155 1336.110 4.280 ;
        RECT 1336.950 0.155 1339.330 4.280 ;
        RECT 1340.170 0.155 1342.550 4.280 ;
        RECT 1343.390 0.155 1345.770 4.280 ;
        RECT 1346.610 0.155 1348.990 4.280 ;
        RECT 1349.830 0.155 1352.210 4.280 ;
        RECT 1353.050 0.155 1355.430 4.280 ;
        RECT 1356.270 0.155 1358.650 4.280 ;
        RECT 1359.490 0.155 1361.870 4.280 ;
        RECT 1362.710 0.155 1365.090 4.280 ;
        RECT 1365.930 0.155 1368.310 4.280 ;
        RECT 1369.150 0.155 1371.530 4.280 ;
        RECT 1372.370 0.155 1374.750 4.280 ;
        RECT 1375.590 0.155 1377.970 4.280 ;
        RECT 1378.810 0.155 1381.190 4.280 ;
        RECT 1382.030 0.155 1387.630 4.280 ;
        RECT 1388.470 0.155 1390.850 4.280 ;
        RECT 1391.690 0.155 1394.070 4.280 ;
        RECT 1394.910 0.155 1397.290 4.280 ;
        RECT 1398.130 0.155 1400.510 4.280 ;
        RECT 1401.350 0.155 1403.730 4.280 ;
        RECT 1404.570 0.155 1406.950 4.280 ;
        RECT 1407.790 0.155 1410.170 4.280 ;
        RECT 1411.010 0.155 1413.390 4.280 ;
        RECT 1414.230 0.155 1416.610 4.280 ;
        RECT 1417.450 0.155 1419.830 4.280 ;
        RECT 1420.670 0.155 1423.050 4.280 ;
        RECT 1423.890 0.155 1426.270 4.280 ;
        RECT 1427.110 0.155 1429.490 4.280 ;
        RECT 1430.330 0.155 1435.930 4.280 ;
        RECT 1436.770 0.155 1439.150 4.280 ;
        RECT 1439.990 0.155 1442.370 4.280 ;
        RECT 1443.210 0.155 1445.590 4.280 ;
        RECT 1446.430 0.155 1448.810 4.280 ;
        RECT 1449.650 0.155 1452.030 4.280 ;
        RECT 1452.870 0.155 1455.250 4.280 ;
        RECT 1456.090 0.155 1458.470 4.280 ;
        RECT 1459.310 0.155 1461.690 4.280 ;
        RECT 1462.530 0.155 1464.910 4.280 ;
        RECT 1465.750 0.155 1468.130 4.280 ;
        RECT 1468.970 0.155 1471.350 4.280 ;
        RECT 1472.190 0.155 1474.570 4.280 ;
        RECT 1475.410 0.155 1477.790 4.280 ;
        RECT 1478.630 0.155 1481.010 4.280 ;
        RECT 1481.850 0.155 1487.450 4.280 ;
        RECT 1488.290 0.155 1490.670 4.280 ;
        RECT 1491.510 0.155 1493.890 4.280 ;
        RECT 1494.730 0.155 1497.110 4.280 ;
        RECT 1497.950 0.155 1500.330 4.280 ;
        RECT 1501.170 0.155 1503.550 4.280 ;
        RECT 1504.390 0.155 1506.770 4.280 ;
        RECT 1507.610 0.155 1509.990 4.280 ;
        RECT 1510.830 0.155 1513.210 4.280 ;
        RECT 1514.050 0.155 1516.430 4.280 ;
        RECT 1517.270 0.155 1519.650 4.280 ;
        RECT 1520.490 0.155 1522.870 4.280 ;
        RECT 1523.710 0.155 1526.090 4.280 ;
        RECT 1526.930 0.155 1529.310 4.280 ;
        RECT 1530.150 0.155 1532.530 4.280 ;
        RECT 1533.370 0.155 1538.970 4.280 ;
        RECT 1539.810 0.155 1542.190 4.280 ;
        RECT 1543.030 0.155 1545.410 4.280 ;
        RECT 1546.250 0.155 1548.630 4.280 ;
        RECT 1549.470 0.155 1551.850 4.280 ;
        RECT 1552.690 0.155 1555.070 4.280 ;
        RECT 1555.910 0.155 1558.290 4.280 ;
        RECT 1559.130 0.155 1561.510 4.280 ;
        RECT 1562.350 0.155 1564.730 4.280 ;
        RECT 1565.570 0.155 1567.950 4.280 ;
        RECT 1568.790 0.155 1571.170 4.280 ;
        RECT 1572.010 0.155 1574.390 4.280 ;
        RECT 1575.230 0.155 1577.610 4.280 ;
        RECT 1578.450 0.155 1580.830 4.280 ;
        RECT 1581.670 0.155 1584.050 4.280 ;
        RECT 1584.890 0.155 1590.490 4.280 ;
        RECT 1591.330 0.155 1593.710 4.280 ;
        RECT 1594.550 0.155 1596.930 4.280 ;
        RECT 1597.770 0.155 1600.150 4.280 ;
        RECT 1600.990 0.155 1603.370 4.280 ;
        RECT 1604.210 0.155 1606.590 4.280 ;
        RECT 1607.430 0.155 1609.810 4.280 ;
        RECT 1610.650 0.155 1613.030 4.280 ;
        RECT 1613.870 0.155 1616.250 4.280 ;
        RECT 1617.090 0.155 1619.470 4.280 ;
        RECT 1620.310 0.155 1622.690 4.280 ;
        RECT 1623.530 0.155 1625.910 4.280 ;
        RECT 1626.750 0.155 1629.130 4.280 ;
        RECT 1629.970 0.155 1632.350 4.280 ;
        RECT 1633.190 0.155 1635.570 4.280 ;
        RECT 1636.410 0.155 1642.010 4.280 ;
        RECT 1642.850 0.155 1645.230 4.280 ;
        RECT 1646.070 0.155 1648.450 4.280 ;
        RECT 1649.290 0.155 1651.670 4.280 ;
        RECT 1652.510 0.155 1654.890 4.280 ;
        RECT 1655.730 0.155 1658.110 4.280 ;
        RECT 1658.950 0.155 1661.330 4.280 ;
        RECT 1662.170 0.155 1664.550 4.280 ;
        RECT 1665.390 0.155 1667.770 4.280 ;
        RECT 1668.610 0.155 1670.990 4.280 ;
        RECT 1671.830 0.155 1674.210 4.280 ;
        RECT 1675.050 0.155 1677.430 4.280 ;
        RECT 1678.270 0.155 1680.650 4.280 ;
        RECT 1681.490 0.155 1683.870 4.280 ;
        RECT 1684.710 0.155 1687.090 4.280 ;
        RECT 1687.930 0.155 1693.530 4.280 ;
        RECT 1694.370 0.155 1696.750 4.280 ;
        RECT 1697.590 0.155 1699.970 4.280 ;
        RECT 1700.810 0.155 1703.190 4.280 ;
        RECT 1704.030 0.155 1706.410 4.280 ;
        RECT 1707.250 0.155 1709.630 4.280 ;
        RECT 1710.470 0.155 1712.850 4.280 ;
        RECT 1713.690 0.155 1716.070 4.280 ;
        RECT 1716.910 0.155 1719.290 4.280 ;
        RECT 1720.130 0.155 1722.510 4.280 ;
        RECT 1723.350 0.155 1725.730 4.280 ;
        RECT 1726.570 0.155 1728.950 4.280 ;
        RECT 1729.790 0.155 1732.170 4.280 ;
        RECT 1733.010 0.155 1735.390 4.280 ;
        RECT 1736.230 0.155 1738.610 4.280 ;
        RECT 1739.450 0.155 1745.050 4.280 ;
        RECT 1745.890 0.155 1748.270 4.280 ;
        RECT 1749.110 0.155 1751.490 4.280 ;
        RECT 1752.330 0.155 1754.710 4.280 ;
        RECT 1755.550 0.155 1757.930 4.280 ;
        RECT 1758.770 0.155 1761.150 4.280 ;
        RECT 1761.990 0.155 1764.370 4.280 ;
        RECT 1765.210 0.155 1767.590 4.280 ;
        RECT 1768.430 0.155 1770.810 4.280 ;
        RECT 1771.650 0.155 1774.030 4.280 ;
        RECT 1774.870 0.155 1777.250 4.280 ;
        RECT 1778.090 0.155 1780.470 4.280 ;
        RECT 1781.310 0.155 1783.690 4.280 ;
        RECT 1784.530 0.155 1786.910 4.280 ;
        RECT 1787.750 0.155 1790.130 4.280 ;
        RECT 1790.970 0.155 1796.570 4.280 ;
        RECT 1797.410 0.155 1799.790 4.280 ;
        RECT 1800.630 0.155 1803.010 4.280 ;
        RECT 1803.850 0.155 1806.230 4.280 ;
        RECT 1807.070 0.155 1809.450 4.280 ;
        RECT 1810.290 0.155 1812.670 4.280 ;
        RECT 1813.510 0.155 1815.890 4.280 ;
        RECT 1816.730 0.155 1819.110 4.280 ;
        RECT 1819.950 0.155 1822.330 4.280 ;
        RECT 1823.170 0.155 1825.550 4.280 ;
        RECT 1826.390 0.155 1828.770 4.280 ;
        RECT 1829.610 0.155 1831.990 4.280 ;
        RECT 1832.830 0.155 1835.210 4.280 ;
        RECT 1836.050 0.155 1838.430 4.280 ;
        RECT 1839.270 0.155 1841.650 4.280 ;
        RECT 1842.490 0.155 1848.090 4.280 ;
        RECT 1848.930 0.155 1851.310 4.280 ;
        RECT 1852.150 0.155 1854.530 4.280 ;
        RECT 1855.370 0.155 1857.750 4.280 ;
        RECT 1858.590 0.155 1860.970 4.280 ;
        RECT 1861.810 0.155 1864.190 4.280 ;
        RECT 1865.030 0.155 1867.410 4.280 ;
        RECT 1868.250 0.155 1870.630 4.280 ;
        RECT 1871.470 0.155 1873.850 4.280 ;
        RECT 1874.690 0.155 1877.070 4.280 ;
        RECT 1877.910 0.155 1880.290 4.280 ;
        RECT 1881.130 0.155 1883.510 4.280 ;
        RECT 1884.350 0.155 1886.730 4.280 ;
        RECT 1887.570 0.155 1889.950 4.280 ;
        RECT 1890.790 0.155 1893.170 4.280 ;
        RECT 1894.010 0.155 1899.610 4.280 ;
        RECT 1900.450 0.155 1902.830 4.280 ;
        RECT 1903.670 0.155 1906.050 4.280 ;
        RECT 1906.890 0.155 1909.270 4.280 ;
        RECT 1910.110 0.155 1912.490 4.280 ;
        RECT 1913.330 0.155 1915.710 4.280 ;
        RECT 1916.550 0.155 1918.930 4.280 ;
        RECT 1919.770 0.155 1922.150 4.280 ;
        RECT 1922.990 0.155 1925.370 4.280 ;
        RECT 1926.210 0.155 1928.590 4.280 ;
        RECT 1929.430 0.155 1931.810 4.280 ;
        RECT 1932.650 0.155 1935.030 4.280 ;
        RECT 1935.870 0.155 1938.250 4.280 ;
        RECT 1939.090 0.155 1941.470 4.280 ;
        RECT 1942.310 0.155 1944.690 4.280 ;
        RECT 1945.530 0.155 1951.130 4.280 ;
        RECT 1951.970 0.155 1954.350 4.280 ;
        RECT 1955.190 0.155 1957.570 4.280 ;
        RECT 1958.410 0.155 1960.790 4.280 ;
        RECT 1961.630 0.155 1964.010 4.280 ;
        RECT 1964.850 0.155 1967.230 4.280 ;
        RECT 1968.070 0.155 1970.450 4.280 ;
        RECT 1971.290 0.155 1973.670 4.280 ;
        RECT 1974.510 0.155 1976.890 4.280 ;
        RECT 1977.730 0.155 1980.110 4.280 ;
        RECT 1980.950 0.155 1983.330 4.280 ;
        RECT 1984.170 0.155 1986.550 4.280 ;
        RECT 1987.390 0.155 1989.770 4.280 ;
        RECT 1990.610 0.155 1992.990 4.280 ;
        RECT 1993.830 0.155 1996.210 4.280 ;
        RECT 1997.050 0.155 2002.650 4.280 ;
        RECT 2003.490 0.155 2005.870 4.280 ;
        RECT 2006.710 0.155 2009.090 4.280 ;
        RECT 2009.930 0.155 2012.310 4.280 ;
        RECT 2013.150 0.155 2015.530 4.280 ;
        RECT 2016.370 0.155 2018.750 4.280 ;
        RECT 2019.590 0.155 2021.970 4.280 ;
        RECT 2022.810 0.155 2025.190 4.280 ;
        RECT 2026.030 0.155 2028.410 4.280 ;
        RECT 2029.250 0.155 2031.630 4.280 ;
        RECT 2032.470 0.155 2034.850 4.280 ;
        RECT 2035.690 0.155 2038.070 4.280 ;
        RECT 2038.910 0.155 2041.290 4.280 ;
        RECT 2042.130 0.155 2044.510 4.280 ;
        RECT 2045.350 0.155 2047.730 4.280 ;
        RECT 2048.570 0.155 2054.170 4.280 ;
        RECT 2055.010 0.155 2057.390 4.280 ;
        RECT 2058.230 0.155 2060.610 4.280 ;
        RECT 2061.450 0.155 2063.830 4.280 ;
        RECT 2064.670 0.155 2067.050 4.280 ;
        RECT 2067.890 0.155 2070.270 4.280 ;
        RECT 2071.110 0.155 2073.490 4.280 ;
        RECT 2074.330 0.155 2076.710 4.280 ;
        RECT 2077.550 0.155 2079.930 4.280 ;
        RECT 2080.770 0.155 2083.150 4.280 ;
        RECT 2083.990 0.155 2086.370 4.280 ;
        RECT 2087.210 0.155 2089.590 4.280 ;
        RECT 2090.430 0.155 2092.810 4.280 ;
        RECT 2093.650 0.155 2096.030 4.280 ;
        RECT 2096.870 0.155 2102.470 4.280 ;
        RECT 2103.310 0.155 2105.690 4.280 ;
        RECT 2106.530 0.155 2108.910 4.280 ;
        RECT 2109.750 0.155 2112.130 4.280 ;
        RECT 2112.970 0.155 2115.350 4.280 ;
        RECT 2116.190 0.155 2118.570 4.280 ;
        RECT 2119.410 0.155 2121.790 4.280 ;
        RECT 2122.630 0.155 2125.010 4.280 ;
        RECT 2125.850 0.155 2128.230 4.280 ;
        RECT 2129.070 0.155 2131.450 4.280 ;
        RECT 2132.290 0.155 2134.670 4.280 ;
        RECT 2135.510 0.155 2137.890 4.280 ;
        RECT 2138.730 0.155 2141.110 4.280 ;
        RECT 2141.950 0.155 2144.330 4.280 ;
        RECT 2145.170 0.155 2147.550 4.280 ;
        RECT 2148.390 0.155 2153.990 4.280 ;
        RECT 2154.830 0.155 2157.210 4.280 ;
        RECT 2158.050 0.155 2160.430 4.280 ;
        RECT 2161.270 0.155 2163.650 4.280 ;
        RECT 2164.490 0.155 2166.870 4.280 ;
        RECT 2167.710 0.155 2170.090 4.280 ;
        RECT 2170.930 0.155 2173.310 4.280 ;
        RECT 2174.150 0.155 2176.530 4.280 ;
        RECT 2177.370 0.155 2179.750 4.280 ;
        RECT 2180.590 0.155 2182.970 4.280 ;
        RECT 2183.810 0.155 2186.190 4.280 ;
        RECT 2187.030 0.155 2189.410 4.280 ;
        RECT 2190.250 0.155 2192.630 4.280 ;
        RECT 2193.470 0.155 2195.850 4.280 ;
        RECT 2196.690 0.155 2199.070 4.280 ;
        RECT 2199.910 0.155 2205.510 4.280 ;
        RECT 2206.350 0.155 2208.730 4.280 ;
        RECT 2209.570 0.155 2211.950 4.280 ;
        RECT 2212.790 0.155 2215.170 4.280 ;
        RECT 2216.010 0.155 2218.390 4.280 ;
        RECT 2219.230 0.155 2221.610 4.280 ;
        RECT 2222.450 0.155 2224.830 4.280 ;
        RECT 2225.670 0.155 2228.050 4.280 ;
        RECT 2228.890 0.155 2231.270 4.280 ;
        RECT 2232.110 0.155 2234.490 4.280 ;
        RECT 2235.330 0.155 2237.710 4.280 ;
        RECT 2238.550 0.155 2240.930 4.280 ;
        RECT 2241.770 0.155 2244.150 4.280 ;
        RECT 2244.990 0.155 2247.370 4.280 ;
        RECT 2248.210 0.155 2250.590 4.280 ;
        RECT 2251.430 0.155 2257.030 4.280 ;
        RECT 2257.870 0.155 2260.250 4.280 ;
        RECT 2261.090 0.155 2263.470 4.280 ;
        RECT 2264.310 0.155 2266.690 4.280 ;
        RECT 2267.530 0.155 2269.910 4.280 ;
        RECT 2270.750 0.155 2273.130 4.280 ;
        RECT 2273.970 0.155 2276.350 4.280 ;
        RECT 2277.190 0.155 2279.570 4.280 ;
        RECT 2280.410 0.155 2282.790 4.280 ;
        RECT 2283.630 0.155 2286.010 4.280 ;
        RECT 2286.850 0.155 2289.230 4.280 ;
        RECT 2290.070 0.155 2292.450 4.280 ;
        RECT 2293.290 0.155 2295.670 4.280 ;
        RECT 2296.510 0.155 2298.890 4.280 ;
        RECT 2299.730 0.155 2302.110 4.280 ;
        RECT 2302.950 0.155 2308.550 4.280 ;
        RECT 2309.390 0.155 2311.770 4.280 ;
        RECT 2312.610 0.155 2314.990 4.280 ;
        RECT 2315.830 0.155 2318.210 4.280 ;
        RECT 2319.050 0.155 2321.430 4.280 ;
        RECT 2322.270 0.155 2324.650 4.280 ;
        RECT 2325.490 0.155 2327.870 4.280 ;
        RECT 2328.710 0.155 2331.090 4.280 ;
        RECT 2331.930 0.155 2334.310 4.280 ;
        RECT 2335.150 0.155 2337.530 4.280 ;
        RECT 2338.370 0.155 2340.750 4.280 ;
        RECT 2341.590 0.155 2343.970 4.280 ;
        RECT 2344.810 0.155 2347.190 4.280 ;
        RECT 2348.030 0.155 2350.410 4.280 ;
        RECT 2351.250 0.155 2353.630 4.280 ;
        RECT 2354.470 0.155 2360.070 4.280 ;
        RECT 2360.910 0.155 2363.290 4.280 ;
        RECT 2364.130 0.155 2366.510 4.280 ;
        RECT 2367.350 0.155 2369.730 4.280 ;
        RECT 2370.570 0.155 2372.950 4.280 ;
        RECT 2373.790 0.155 2376.170 4.280 ;
        RECT 2377.010 0.155 2379.390 4.280 ;
        RECT 2380.230 0.155 2382.610 4.280 ;
        RECT 2383.450 0.155 2385.830 4.280 ;
        RECT 2386.670 0.155 2389.050 4.280 ;
        RECT 2389.890 0.155 2392.270 4.280 ;
        RECT 2393.110 0.155 2395.490 4.280 ;
        RECT 2396.330 0.155 2398.710 4.280 ;
        RECT 2399.550 0.155 2401.930 4.280 ;
        RECT 2402.770 0.155 2405.150 4.280 ;
        RECT 2405.990 0.155 2411.590 4.280 ;
        RECT 2412.430 0.155 2414.810 4.280 ;
        RECT 2415.650 0.155 2418.030 4.280 ;
        RECT 2418.870 0.155 2421.250 4.280 ;
        RECT 2422.090 0.155 2424.470 4.280 ;
        RECT 2425.310 0.155 2427.690 4.280 ;
        RECT 2428.530 0.155 2430.910 4.280 ;
        RECT 2431.750 0.155 2434.130 4.280 ;
        RECT 2434.970 0.155 2437.350 4.280 ;
        RECT 2438.190 0.155 2440.570 4.280 ;
        RECT 2441.410 0.155 2443.790 4.280 ;
        RECT 2444.630 0.155 2447.010 4.280 ;
        RECT 2447.850 0.155 2450.230 4.280 ;
        RECT 2451.070 0.155 2453.450 4.280 ;
        RECT 2454.290 0.155 2456.670 4.280 ;
        RECT 2457.510 0.155 2463.110 4.280 ;
        RECT 2463.950 0.155 2466.330 4.280 ;
        RECT 2467.170 0.155 2469.550 4.280 ;
        RECT 2470.390 0.155 2472.770 4.280 ;
        RECT 2473.610 0.155 2475.990 4.280 ;
        RECT 2476.830 0.155 2479.210 4.280 ;
        RECT 2480.050 0.155 2482.430 4.280 ;
        RECT 2483.270 0.155 2485.650 4.280 ;
        RECT 2486.490 0.155 2488.870 4.280 ;
        RECT 2489.710 0.155 2492.090 4.280 ;
        RECT 2492.930 0.155 2495.310 4.280 ;
        RECT 2496.150 0.155 2498.530 4.280 ;
      LAYER met3 ;
        RECT 4.400 2498.640 2498.195 2499.505 ;
        RECT 4.000 2496.640 2498.195 2498.640 ;
        RECT 4.400 2495.240 2495.600 2496.640 ;
        RECT 4.000 2493.240 2498.195 2495.240 ;
        RECT 4.400 2491.840 2495.600 2493.240 ;
        RECT 4.000 2489.840 2498.195 2491.840 ;
        RECT 4.000 2488.440 2495.600 2489.840 ;
        RECT 4.000 2486.440 2498.195 2488.440 ;
        RECT 4.400 2485.040 2495.600 2486.440 ;
        RECT 4.000 2483.040 2498.195 2485.040 ;
        RECT 4.400 2481.640 2495.600 2483.040 ;
        RECT 4.000 2479.640 2498.195 2481.640 ;
        RECT 4.400 2478.240 2495.600 2479.640 ;
        RECT 4.000 2476.240 2498.195 2478.240 ;
        RECT 4.400 2474.840 2495.600 2476.240 ;
        RECT 4.000 2472.840 2498.195 2474.840 ;
        RECT 4.400 2471.440 2495.600 2472.840 ;
        RECT 4.000 2469.440 2498.195 2471.440 ;
        RECT 4.400 2468.040 2495.600 2469.440 ;
        RECT 4.000 2466.040 2498.195 2468.040 ;
        RECT 4.400 2464.640 2495.600 2466.040 ;
        RECT 4.000 2462.640 2498.195 2464.640 ;
        RECT 4.400 2461.240 2495.600 2462.640 ;
        RECT 4.000 2459.240 2498.195 2461.240 ;
        RECT 4.400 2457.840 2495.600 2459.240 ;
        RECT 4.000 2455.840 2498.195 2457.840 ;
        RECT 4.400 2454.440 2495.600 2455.840 ;
        RECT 4.000 2452.440 2498.195 2454.440 ;
        RECT 4.400 2451.040 2495.600 2452.440 ;
        RECT 4.000 2449.040 2498.195 2451.040 ;
        RECT 4.400 2447.640 2498.195 2449.040 ;
        RECT 4.000 2445.640 2498.195 2447.640 ;
        RECT 4.400 2444.240 2495.600 2445.640 ;
        RECT 4.000 2442.240 2498.195 2444.240 ;
        RECT 4.400 2440.840 2495.600 2442.240 ;
        RECT 4.000 2438.840 2498.195 2440.840 ;
        RECT 4.400 2437.440 2495.600 2438.840 ;
        RECT 4.000 2435.440 2498.195 2437.440 ;
        RECT 4.000 2434.040 2495.600 2435.440 ;
        RECT 4.000 2432.040 2498.195 2434.040 ;
        RECT 4.400 2430.640 2495.600 2432.040 ;
        RECT 4.000 2428.640 2498.195 2430.640 ;
        RECT 4.400 2427.240 2495.600 2428.640 ;
        RECT 4.000 2425.240 2498.195 2427.240 ;
        RECT 4.400 2423.840 2495.600 2425.240 ;
        RECT 4.000 2421.840 2498.195 2423.840 ;
        RECT 4.400 2420.440 2495.600 2421.840 ;
        RECT 4.000 2418.440 2498.195 2420.440 ;
        RECT 4.400 2417.040 2495.600 2418.440 ;
        RECT 4.000 2415.040 2498.195 2417.040 ;
        RECT 4.400 2413.640 2495.600 2415.040 ;
        RECT 4.000 2411.640 2498.195 2413.640 ;
        RECT 4.400 2410.240 2495.600 2411.640 ;
        RECT 4.000 2408.240 2498.195 2410.240 ;
        RECT 4.400 2406.840 2495.600 2408.240 ;
        RECT 4.000 2404.840 2498.195 2406.840 ;
        RECT 4.400 2403.440 2495.600 2404.840 ;
        RECT 4.000 2401.440 2498.195 2403.440 ;
        RECT 4.400 2400.040 2495.600 2401.440 ;
        RECT 4.000 2398.040 2498.195 2400.040 ;
        RECT 4.400 2396.640 2495.600 2398.040 ;
        RECT 4.000 2394.640 2498.195 2396.640 ;
        RECT 4.400 2393.240 2498.195 2394.640 ;
        RECT 4.000 2391.240 2498.195 2393.240 ;
        RECT 4.400 2389.840 2495.600 2391.240 ;
        RECT 4.000 2387.840 2498.195 2389.840 ;
        RECT 4.400 2386.440 2495.600 2387.840 ;
        RECT 4.000 2384.440 2498.195 2386.440 ;
        RECT 4.400 2383.040 2495.600 2384.440 ;
        RECT 4.000 2381.040 2498.195 2383.040 ;
        RECT 4.000 2379.640 2495.600 2381.040 ;
        RECT 4.000 2377.640 2498.195 2379.640 ;
        RECT 4.400 2376.240 2495.600 2377.640 ;
        RECT 4.000 2374.240 2498.195 2376.240 ;
        RECT 4.400 2372.840 2495.600 2374.240 ;
        RECT 4.000 2370.840 2498.195 2372.840 ;
        RECT 4.400 2369.440 2495.600 2370.840 ;
        RECT 4.000 2367.440 2498.195 2369.440 ;
        RECT 4.400 2366.040 2495.600 2367.440 ;
        RECT 4.000 2364.040 2498.195 2366.040 ;
        RECT 4.400 2362.640 2495.600 2364.040 ;
        RECT 4.000 2360.640 2498.195 2362.640 ;
        RECT 4.400 2359.240 2495.600 2360.640 ;
        RECT 4.000 2357.240 2498.195 2359.240 ;
        RECT 4.400 2355.840 2495.600 2357.240 ;
        RECT 4.000 2353.840 2498.195 2355.840 ;
        RECT 4.400 2352.440 2495.600 2353.840 ;
        RECT 4.000 2350.440 2498.195 2352.440 ;
        RECT 4.400 2349.040 2495.600 2350.440 ;
        RECT 4.000 2347.040 2498.195 2349.040 ;
        RECT 4.400 2345.640 2495.600 2347.040 ;
        RECT 4.000 2343.640 2498.195 2345.640 ;
        RECT 4.400 2342.240 2495.600 2343.640 ;
        RECT 4.000 2340.240 2498.195 2342.240 ;
        RECT 4.400 2338.840 2498.195 2340.240 ;
        RECT 4.000 2336.840 2498.195 2338.840 ;
        RECT 4.400 2335.440 2495.600 2336.840 ;
        RECT 4.000 2333.440 2498.195 2335.440 ;
        RECT 4.400 2332.040 2495.600 2333.440 ;
        RECT 4.000 2330.040 2498.195 2332.040 ;
        RECT 4.400 2328.640 2495.600 2330.040 ;
        RECT 4.000 2326.640 2498.195 2328.640 ;
        RECT 4.000 2325.240 2495.600 2326.640 ;
        RECT 4.000 2323.240 2498.195 2325.240 ;
        RECT 4.400 2321.840 2495.600 2323.240 ;
        RECT 4.000 2319.840 2498.195 2321.840 ;
        RECT 4.400 2318.440 2495.600 2319.840 ;
        RECT 4.000 2316.440 2498.195 2318.440 ;
        RECT 4.400 2315.040 2495.600 2316.440 ;
        RECT 4.000 2313.040 2498.195 2315.040 ;
        RECT 4.400 2311.640 2495.600 2313.040 ;
        RECT 4.000 2309.640 2498.195 2311.640 ;
        RECT 4.400 2308.240 2495.600 2309.640 ;
        RECT 4.000 2306.240 2498.195 2308.240 ;
        RECT 4.400 2304.840 2495.600 2306.240 ;
        RECT 4.000 2302.840 2498.195 2304.840 ;
        RECT 4.400 2301.440 2495.600 2302.840 ;
        RECT 4.000 2299.440 2498.195 2301.440 ;
        RECT 4.400 2298.040 2495.600 2299.440 ;
        RECT 4.000 2296.040 2498.195 2298.040 ;
        RECT 4.400 2294.640 2495.600 2296.040 ;
        RECT 4.000 2292.640 2498.195 2294.640 ;
        RECT 4.400 2291.240 2495.600 2292.640 ;
        RECT 4.000 2289.240 2498.195 2291.240 ;
        RECT 4.400 2287.840 2495.600 2289.240 ;
        RECT 4.000 2285.840 2498.195 2287.840 ;
        RECT 4.400 2284.440 2498.195 2285.840 ;
        RECT 4.000 2282.440 2498.195 2284.440 ;
        RECT 4.400 2281.040 2495.600 2282.440 ;
        RECT 4.000 2279.040 2498.195 2281.040 ;
        RECT 4.400 2277.640 2495.600 2279.040 ;
        RECT 4.000 2275.640 2498.195 2277.640 ;
        RECT 4.400 2274.240 2495.600 2275.640 ;
        RECT 4.000 2272.240 2498.195 2274.240 ;
        RECT 4.000 2270.840 2495.600 2272.240 ;
        RECT 4.000 2268.840 2498.195 2270.840 ;
        RECT 4.400 2267.440 2495.600 2268.840 ;
        RECT 4.000 2265.440 2498.195 2267.440 ;
        RECT 4.400 2264.040 2495.600 2265.440 ;
        RECT 4.000 2262.040 2498.195 2264.040 ;
        RECT 4.400 2260.640 2495.600 2262.040 ;
        RECT 4.000 2258.640 2498.195 2260.640 ;
        RECT 4.400 2257.240 2495.600 2258.640 ;
        RECT 4.000 2255.240 2498.195 2257.240 ;
        RECT 4.400 2253.840 2495.600 2255.240 ;
        RECT 4.000 2251.840 2498.195 2253.840 ;
        RECT 4.400 2250.440 2495.600 2251.840 ;
        RECT 4.000 2248.440 2498.195 2250.440 ;
        RECT 4.400 2247.040 2495.600 2248.440 ;
        RECT 4.000 2245.040 2498.195 2247.040 ;
        RECT 4.400 2243.640 2495.600 2245.040 ;
        RECT 4.000 2241.640 2498.195 2243.640 ;
        RECT 4.400 2240.240 2495.600 2241.640 ;
        RECT 4.000 2238.240 2498.195 2240.240 ;
        RECT 4.400 2236.840 2495.600 2238.240 ;
        RECT 4.000 2234.840 2498.195 2236.840 ;
        RECT 4.400 2233.440 2495.600 2234.840 ;
        RECT 4.000 2231.440 2498.195 2233.440 ;
        RECT 4.400 2230.040 2498.195 2231.440 ;
        RECT 4.000 2228.040 2498.195 2230.040 ;
        RECT 4.400 2226.640 2495.600 2228.040 ;
        RECT 4.000 2224.640 2498.195 2226.640 ;
        RECT 4.400 2223.240 2495.600 2224.640 ;
        RECT 4.000 2221.240 2498.195 2223.240 ;
        RECT 4.400 2219.840 2495.600 2221.240 ;
        RECT 4.000 2217.840 2498.195 2219.840 ;
        RECT 4.000 2216.440 2495.600 2217.840 ;
        RECT 4.000 2214.440 2498.195 2216.440 ;
        RECT 4.400 2213.040 2495.600 2214.440 ;
        RECT 4.000 2211.040 2498.195 2213.040 ;
        RECT 4.400 2209.640 2495.600 2211.040 ;
        RECT 4.000 2207.640 2498.195 2209.640 ;
        RECT 4.400 2206.240 2495.600 2207.640 ;
        RECT 4.000 2204.240 2498.195 2206.240 ;
        RECT 4.400 2202.840 2495.600 2204.240 ;
        RECT 4.000 2200.840 2498.195 2202.840 ;
        RECT 4.400 2199.440 2495.600 2200.840 ;
        RECT 4.000 2197.440 2498.195 2199.440 ;
        RECT 4.400 2196.040 2495.600 2197.440 ;
        RECT 4.000 2194.040 2498.195 2196.040 ;
        RECT 4.400 2192.640 2495.600 2194.040 ;
        RECT 4.000 2190.640 2498.195 2192.640 ;
        RECT 4.400 2189.240 2495.600 2190.640 ;
        RECT 4.000 2187.240 2498.195 2189.240 ;
        RECT 4.400 2185.840 2495.600 2187.240 ;
        RECT 4.000 2183.840 2498.195 2185.840 ;
        RECT 4.400 2182.440 2495.600 2183.840 ;
        RECT 4.000 2180.440 2498.195 2182.440 ;
        RECT 4.400 2179.040 2495.600 2180.440 ;
        RECT 4.000 2177.040 2498.195 2179.040 ;
        RECT 4.400 2175.640 2498.195 2177.040 ;
        RECT 4.000 2173.640 2498.195 2175.640 ;
        RECT 4.400 2172.240 2495.600 2173.640 ;
        RECT 4.000 2170.240 2498.195 2172.240 ;
        RECT 4.400 2168.840 2495.600 2170.240 ;
        RECT 4.000 2166.840 2498.195 2168.840 ;
        RECT 4.000 2165.440 2495.600 2166.840 ;
        RECT 4.000 2163.440 2498.195 2165.440 ;
        RECT 4.400 2162.040 2495.600 2163.440 ;
        RECT 4.000 2160.040 2498.195 2162.040 ;
        RECT 4.400 2158.640 2495.600 2160.040 ;
        RECT 4.000 2156.640 2498.195 2158.640 ;
        RECT 4.400 2155.240 2495.600 2156.640 ;
        RECT 4.000 2153.240 2498.195 2155.240 ;
        RECT 4.400 2151.840 2495.600 2153.240 ;
        RECT 4.000 2149.840 2498.195 2151.840 ;
        RECT 4.400 2148.440 2495.600 2149.840 ;
        RECT 4.000 2146.440 2498.195 2148.440 ;
        RECT 4.400 2145.040 2495.600 2146.440 ;
        RECT 4.000 2143.040 2498.195 2145.040 ;
        RECT 4.400 2141.640 2495.600 2143.040 ;
        RECT 4.000 2139.640 2498.195 2141.640 ;
        RECT 4.400 2138.240 2495.600 2139.640 ;
        RECT 4.000 2136.240 2498.195 2138.240 ;
        RECT 4.400 2134.840 2495.600 2136.240 ;
        RECT 4.000 2132.840 2498.195 2134.840 ;
        RECT 4.400 2131.440 2495.600 2132.840 ;
        RECT 4.000 2129.440 2498.195 2131.440 ;
        RECT 4.400 2128.040 2495.600 2129.440 ;
        RECT 4.000 2126.040 2498.195 2128.040 ;
        RECT 4.400 2124.640 2495.600 2126.040 ;
        RECT 4.000 2122.640 2498.195 2124.640 ;
        RECT 4.400 2121.240 2498.195 2122.640 ;
        RECT 4.000 2119.240 2498.195 2121.240 ;
        RECT 4.400 2117.840 2495.600 2119.240 ;
        RECT 4.000 2115.840 2498.195 2117.840 ;
        RECT 4.400 2114.440 2495.600 2115.840 ;
        RECT 4.000 2112.440 2498.195 2114.440 ;
        RECT 4.000 2111.040 2495.600 2112.440 ;
        RECT 4.000 2109.040 2498.195 2111.040 ;
        RECT 4.400 2107.640 2495.600 2109.040 ;
        RECT 4.000 2105.640 2498.195 2107.640 ;
        RECT 4.400 2104.240 2495.600 2105.640 ;
        RECT 4.000 2102.240 2498.195 2104.240 ;
        RECT 4.400 2100.840 2495.600 2102.240 ;
        RECT 4.000 2098.840 2498.195 2100.840 ;
        RECT 4.400 2097.440 2495.600 2098.840 ;
        RECT 4.000 2095.440 2498.195 2097.440 ;
        RECT 4.400 2094.040 2495.600 2095.440 ;
        RECT 4.000 2092.040 2498.195 2094.040 ;
        RECT 4.400 2090.640 2495.600 2092.040 ;
        RECT 4.000 2088.640 2498.195 2090.640 ;
        RECT 4.400 2087.240 2495.600 2088.640 ;
        RECT 4.000 2085.240 2498.195 2087.240 ;
        RECT 4.400 2083.840 2495.600 2085.240 ;
        RECT 4.000 2081.840 2498.195 2083.840 ;
        RECT 4.400 2080.440 2495.600 2081.840 ;
        RECT 4.000 2078.440 2498.195 2080.440 ;
        RECT 4.400 2077.040 2495.600 2078.440 ;
        RECT 4.000 2075.040 2498.195 2077.040 ;
        RECT 4.400 2073.640 2495.600 2075.040 ;
        RECT 4.000 2071.640 2498.195 2073.640 ;
        RECT 4.400 2070.240 2495.600 2071.640 ;
        RECT 4.000 2068.240 2498.195 2070.240 ;
        RECT 4.400 2066.840 2498.195 2068.240 ;
        RECT 4.000 2064.840 2498.195 2066.840 ;
        RECT 4.400 2063.440 2495.600 2064.840 ;
        RECT 4.000 2061.440 2498.195 2063.440 ;
        RECT 4.400 2060.040 2495.600 2061.440 ;
        RECT 4.000 2058.040 2498.195 2060.040 ;
        RECT 4.000 2056.640 2495.600 2058.040 ;
        RECT 4.000 2054.640 2498.195 2056.640 ;
        RECT 4.400 2053.240 2495.600 2054.640 ;
        RECT 4.000 2051.240 2498.195 2053.240 ;
        RECT 4.400 2049.840 2495.600 2051.240 ;
        RECT 4.000 2047.840 2498.195 2049.840 ;
        RECT 4.400 2046.440 2495.600 2047.840 ;
        RECT 4.000 2044.440 2498.195 2046.440 ;
        RECT 4.400 2043.040 2495.600 2044.440 ;
        RECT 4.000 2041.040 2498.195 2043.040 ;
        RECT 4.400 2039.640 2495.600 2041.040 ;
        RECT 4.000 2037.640 2498.195 2039.640 ;
        RECT 4.400 2036.240 2495.600 2037.640 ;
        RECT 4.000 2034.240 2498.195 2036.240 ;
        RECT 4.400 2032.840 2495.600 2034.240 ;
        RECT 4.000 2030.840 2498.195 2032.840 ;
        RECT 4.400 2029.440 2495.600 2030.840 ;
        RECT 4.000 2027.440 2498.195 2029.440 ;
        RECT 4.400 2026.040 2495.600 2027.440 ;
        RECT 4.000 2024.040 2498.195 2026.040 ;
        RECT 4.400 2022.640 2495.600 2024.040 ;
        RECT 4.000 2020.640 2498.195 2022.640 ;
        RECT 4.400 2019.240 2495.600 2020.640 ;
        RECT 4.000 2017.240 2498.195 2019.240 ;
        RECT 4.400 2015.840 2495.600 2017.240 ;
        RECT 4.000 2013.840 2498.195 2015.840 ;
        RECT 4.400 2012.440 2498.195 2013.840 ;
        RECT 4.000 2010.440 2498.195 2012.440 ;
        RECT 4.400 2009.040 2495.600 2010.440 ;
        RECT 4.000 2007.040 2498.195 2009.040 ;
        RECT 4.400 2005.640 2495.600 2007.040 ;
        RECT 4.000 2003.640 2498.195 2005.640 ;
        RECT 4.000 2002.240 2495.600 2003.640 ;
        RECT 4.000 2000.240 2498.195 2002.240 ;
        RECT 4.400 1998.840 2495.600 2000.240 ;
        RECT 4.000 1996.840 2498.195 1998.840 ;
        RECT 4.400 1995.440 2495.600 1996.840 ;
        RECT 4.000 1993.440 2498.195 1995.440 ;
        RECT 4.400 1992.040 2495.600 1993.440 ;
        RECT 4.000 1990.040 2498.195 1992.040 ;
        RECT 4.400 1988.640 2495.600 1990.040 ;
        RECT 4.000 1986.640 2498.195 1988.640 ;
        RECT 4.400 1985.240 2495.600 1986.640 ;
        RECT 4.000 1983.240 2498.195 1985.240 ;
        RECT 4.400 1981.840 2495.600 1983.240 ;
        RECT 4.000 1979.840 2498.195 1981.840 ;
        RECT 4.400 1978.440 2495.600 1979.840 ;
        RECT 4.000 1976.440 2498.195 1978.440 ;
        RECT 4.400 1975.040 2495.600 1976.440 ;
        RECT 4.000 1973.040 2498.195 1975.040 ;
        RECT 4.400 1971.640 2495.600 1973.040 ;
        RECT 4.000 1969.640 2498.195 1971.640 ;
        RECT 4.400 1968.240 2495.600 1969.640 ;
        RECT 4.000 1966.240 2498.195 1968.240 ;
        RECT 4.400 1964.840 2495.600 1966.240 ;
        RECT 4.000 1962.840 2498.195 1964.840 ;
        RECT 4.400 1961.440 2495.600 1962.840 ;
        RECT 4.000 1959.440 2498.195 1961.440 ;
        RECT 4.400 1958.040 2498.195 1959.440 ;
        RECT 4.000 1956.040 2498.195 1958.040 ;
        RECT 4.400 1954.640 2495.600 1956.040 ;
        RECT 4.000 1952.640 2498.195 1954.640 ;
        RECT 4.400 1951.240 2495.600 1952.640 ;
        RECT 4.000 1949.240 2498.195 1951.240 ;
        RECT 4.000 1947.840 2495.600 1949.240 ;
        RECT 4.000 1945.840 2498.195 1947.840 ;
        RECT 4.400 1944.440 2495.600 1945.840 ;
        RECT 4.000 1942.440 2498.195 1944.440 ;
        RECT 4.400 1941.040 2495.600 1942.440 ;
        RECT 4.000 1939.040 2498.195 1941.040 ;
        RECT 4.400 1937.640 2495.600 1939.040 ;
        RECT 4.000 1935.640 2498.195 1937.640 ;
        RECT 4.400 1934.240 2495.600 1935.640 ;
        RECT 4.000 1932.240 2498.195 1934.240 ;
        RECT 4.400 1930.840 2495.600 1932.240 ;
        RECT 4.000 1928.840 2498.195 1930.840 ;
        RECT 4.400 1927.440 2495.600 1928.840 ;
        RECT 4.000 1925.440 2498.195 1927.440 ;
        RECT 4.400 1924.040 2495.600 1925.440 ;
        RECT 4.000 1922.040 2498.195 1924.040 ;
        RECT 4.400 1920.640 2495.600 1922.040 ;
        RECT 4.000 1918.640 2498.195 1920.640 ;
        RECT 4.400 1917.240 2495.600 1918.640 ;
        RECT 4.000 1915.240 2498.195 1917.240 ;
        RECT 4.400 1913.840 2495.600 1915.240 ;
        RECT 4.000 1911.840 2498.195 1913.840 ;
        RECT 4.400 1910.440 2495.600 1911.840 ;
        RECT 4.000 1908.440 2498.195 1910.440 ;
        RECT 4.400 1907.040 2495.600 1908.440 ;
        RECT 4.000 1905.040 2498.195 1907.040 ;
        RECT 4.400 1903.640 2498.195 1905.040 ;
        RECT 4.000 1901.640 2498.195 1903.640 ;
        RECT 4.400 1900.240 2495.600 1901.640 ;
        RECT 4.000 1898.240 2498.195 1900.240 ;
        RECT 4.400 1896.840 2495.600 1898.240 ;
        RECT 4.000 1894.840 2498.195 1896.840 ;
        RECT 4.000 1893.440 2495.600 1894.840 ;
        RECT 4.000 1891.440 2498.195 1893.440 ;
        RECT 4.400 1890.040 2495.600 1891.440 ;
        RECT 4.000 1888.040 2498.195 1890.040 ;
        RECT 4.400 1886.640 2495.600 1888.040 ;
        RECT 4.000 1884.640 2498.195 1886.640 ;
        RECT 4.400 1883.240 2495.600 1884.640 ;
        RECT 4.000 1881.240 2498.195 1883.240 ;
        RECT 4.400 1879.840 2495.600 1881.240 ;
        RECT 4.000 1877.840 2498.195 1879.840 ;
        RECT 4.400 1876.440 2495.600 1877.840 ;
        RECT 4.000 1874.440 2498.195 1876.440 ;
        RECT 4.400 1873.040 2495.600 1874.440 ;
        RECT 4.000 1871.040 2498.195 1873.040 ;
        RECT 4.400 1869.640 2495.600 1871.040 ;
        RECT 4.000 1867.640 2498.195 1869.640 ;
        RECT 4.400 1866.240 2495.600 1867.640 ;
        RECT 4.000 1864.240 2498.195 1866.240 ;
        RECT 4.400 1862.840 2495.600 1864.240 ;
        RECT 4.000 1860.840 2498.195 1862.840 ;
        RECT 4.400 1859.440 2495.600 1860.840 ;
        RECT 4.000 1857.440 2498.195 1859.440 ;
        RECT 4.400 1856.040 2495.600 1857.440 ;
        RECT 4.000 1854.040 2498.195 1856.040 ;
        RECT 4.400 1852.640 2495.600 1854.040 ;
        RECT 4.000 1850.640 2498.195 1852.640 ;
        RECT 4.400 1849.240 2498.195 1850.640 ;
        RECT 4.000 1847.240 2498.195 1849.240 ;
        RECT 4.400 1845.840 2495.600 1847.240 ;
        RECT 4.000 1843.840 2498.195 1845.840 ;
        RECT 4.400 1842.440 2495.600 1843.840 ;
        RECT 4.000 1840.440 2498.195 1842.440 ;
        RECT 4.000 1839.040 2495.600 1840.440 ;
        RECT 4.000 1837.040 2498.195 1839.040 ;
        RECT 4.400 1835.640 2495.600 1837.040 ;
        RECT 4.000 1833.640 2498.195 1835.640 ;
        RECT 4.400 1832.240 2495.600 1833.640 ;
        RECT 4.000 1830.240 2498.195 1832.240 ;
        RECT 4.400 1828.840 2495.600 1830.240 ;
        RECT 4.000 1826.840 2498.195 1828.840 ;
        RECT 4.400 1825.440 2495.600 1826.840 ;
        RECT 4.000 1823.440 2498.195 1825.440 ;
        RECT 4.400 1822.040 2495.600 1823.440 ;
        RECT 4.000 1820.040 2498.195 1822.040 ;
        RECT 4.400 1818.640 2495.600 1820.040 ;
        RECT 4.000 1816.640 2498.195 1818.640 ;
        RECT 4.400 1815.240 2495.600 1816.640 ;
        RECT 4.000 1813.240 2498.195 1815.240 ;
        RECT 4.400 1811.840 2495.600 1813.240 ;
        RECT 4.000 1809.840 2498.195 1811.840 ;
        RECT 4.400 1808.440 2495.600 1809.840 ;
        RECT 4.000 1806.440 2498.195 1808.440 ;
        RECT 4.400 1805.040 2495.600 1806.440 ;
        RECT 4.000 1803.040 2498.195 1805.040 ;
        RECT 4.400 1801.640 2495.600 1803.040 ;
        RECT 4.000 1799.640 2498.195 1801.640 ;
        RECT 4.400 1798.240 2495.600 1799.640 ;
        RECT 4.000 1796.240 2498.195 1798.240 ;
        RECT 4.400 1794.840 2498.195 1796.240 ;
        RECT 4.000 1792.840 2498.195 1794.840 ;
        RECT 4.400 1791.440 2495.600 1792.840 ;
        RECT 4.000 1789.440 2498.195 1791.440 ;
        RECT 4.400 1788.040 2495.600 1789.440 ;
        RECT 4.000 1786.040 2498.195 1788.040 ;
        RECT 4.000 1784.640 2495.600 1786.040 ;
        RECT 4.000 1782.640 2498.195 1784.640 ;
        RECT 4.400 1781.240 2495.600 1782.640 ;
        RECT 4.000 1779.240 2498.195 1781.240 ;
        RECT 4.400 1777.840 2495.600 1779.240 ;
        RECT 4.000 1775.840 2498.195 1777.840 ;
        RECT 4.400 1774.440 2495.600 1775.840 ;
        RECT 4.000 1772.440 2498.195 1774.440 ;
        RECT 4.400 1771.040 2495.600 1772.440 ;
        RECT 4.000 1769.040 2498.195 1771.040 ;
        RECT 4.400 1767.640 2495.600 1769.040 ;
        RECT 4.000 1765.640 2498.195 1767.640 ;
        RECT 4.400 1764.240 2495.600 1765.640 ;
        RECT 4.000 1762.240 2498.195 1764.240 ;
        RECT 4.400 1760.840 2495.600 1762.240 ;
        RECT 4.000 1758.840 2498.195 1760.840 ;
        RECT 4.400 1757.440 2495.600 1758.840 ;
        RECT 4.000 1755.440 2498.195 1757.440 ;
        RECT 4.400 1754.040 2495.600 1755.440 ;
        RECT 4.000 1752.040 2498.195 1754.040 ;
        RECT 4.400 1750.640 2495.600 1752.040 ;
        RECT 4.000 1748.640 2498.195 1750.640 ;
        RECT 4.400 1747.240 2495.600 1748.640 ;
        RECT 4.000 1745.240 2498.195 1747.240 ;
        RECT 4.400 1743.840 2498.195 1745.240 ;
        RECT 4.000 1741.840 2498.195 1743.840 ;
        RECT 4.400 1740.440 2495.600 1741.840 ;
        RECT 4.000 1738.440 2498.195 1740.440 ;
        RECT 4.400 1737.040 2495.600 1738.440 ;
        RECT 4.000 1735.040 2498.195 1737.040 ;
        RECT 4.400 1733.640 2495.600 1735.040 ;
        RECT 4.000 1731.640 2498.195 1733.640 ;
        RECT 4.000 1730.240 2495.600 1731.640 ;
        RECT 4.000 1728.240 2498.195 1730.240 ;
        RECT 4.400 1726.840 2495.600 1728.240 ;
        RECT 4.000 1724.840 2498.195 1726.840 ;
        RECT 4.400 1723.440 2495.600 1724.840 ;
        RECT 4.000 1721.440 2498.195 1723.440 ;
        RECT 4.400 1720.040 2495.600 1721.440 ;
        RECT 4.000 1718.040 2498.195 1720.040 ;
        RECT 4.400 1716.640 2495.600 1718.040 ;
        RECT 4.000 1714.640 2498.195 1716.640 ;
        RECT 4.400 1713.240 2495.600 1714.640 ;
        RECT 4.000 1711.240 2498.195 1713.240 ;
        RECT 4.400 1709.840 2495.600 1711.240 ;
        RECT 4.000 1707.840 2498.195 1709.840 ;
        RECT 4.400 1706.440 2495.600 1707.840 ;
        RECT 4.000 1704.440 2498.195 1706.440 ;
        RECT 4.400 1703.040 2495.600 1704.440 ;
        RECT 4.000 1701.040 2498.195 1703.040 ;
        RECT 4.400 1699.640 2495.600 1701.040 ;
        RECT 4.000 1697.640 2498.195 1699.640 ;
        RECT 4.400 1696.240 2495.600 1697.640 ;
        RECT 4.000 1694.240 2498.195 1696.240 ;
        RECT 4.400 1692.840 2495.600 1694.240 ;
        RECT 4.000 1690.840 2498.195 1692.840 ;
        RECT 4.400 1689.440 2498.195 1690.840 ;
        RECT 4.000 1687.440 2498.195 1689.440 ;
        RECT 4.400 1686.040 2495.600 1687.440 ;
        RECT 4.000 1684.040 2498.195 1686.040 ;
        RECT 4.400 1682.640 2495.600 1684.040 ;
        RECT 4.000 1680.640 2498.195 1682.640 ;
        RECT 4.400 1679.240 2495.600 1680.640 ;
        RECT 4.000 1677.240 2498.195 1679.240 ;
        RECT 4.000 1675.840 2495.600 1677.240 ;
        RECT 4.000 1673.840 2498.195 1675.840 ;
        RECT 4.400 1672.440 2495.600 1673.840 ;
        RECT 4.000 1670.440 2498.195 1672.440 ;
        RECT 4.400 1669.040 2495.600 1670.440 ;
        RECT 4.000 1667.040 2498.195 1669.040 ;
        RECT 4.400 1665.640 2495.600 1667.040 ;
        RECT 4.000 1663.640 2498.195 1665.640 ;
        RECT 4.400 1662.240 2495.600 1663.640 ;
        RECT 4.000 1660.240 2498.195 1662.240 ;
        RECT 4.400 1658.840 2495.600 1660.240 ;
        RECT 4.000 1656.840 2498.195 1658.840 ;
        RECT 4.400 1655.440 2495.600 1656.840 ;
        RECT 4.000 1653.440 2498.195 1655.440 ;
        RECT 4.400 1652.040 2495.600 1653.440 ;
        RECT 4.000 1650.040 2498.195 1652.040 ;
        RECT 4.400 1648.640 2495.600 1650.040 ;
        RECT 4.000 1646.640 2498.195 1648.640 ;
        RECT 4.400 1645.240 2495.600 1646.640 ;
        RECT 4.000 1643.240 2498.195 1645.240 ;
        RECT 4.400 1641.840 2495.600 1643.240 ;
        RECT 4.000 1639.840 2498.195 1641.840 ;
        RECT 4.400 1638.440 2495.600 1639.840 ;
        RECT 4.000 1636.440 2498.195 1638.440 ;
        RECT 4.400 1635.040 2498.195 1636.440 ;
        RECT 4.000 1633.040 2498.195 1635.040 ;
        RECT 4.400 1631.640 2495.600 1633.040 ;
        RECT 4.000 1629.640 2498.195 1631.640 ;
        RECT 4.400 1628.240 2495.600 1629.640 ;
        RECT 4.000 1626.240 2498.195 1628.240 ;
        RECT 4.400 1624.840 2495.600 1626.240 ;
        RECT 4.000 1622.840 2498.195 1624.840 ;
        RECT 4.000 1621.440 2495.600 1622.840 ;
        RECT 4.000 1619.440 2498.195 1621.440 ;
        RECT 4.400 1618.040 2495.600 1619.440 ;
        RECT 4.000 1616.040 2498.195 1618.040 ;
        RECT 4.400 1614.640 2495.600 1616.040 ;
        RECT 4.000 1612.640 2498.195 1614.640 ;
        RECT 4.400 1611.240 2495.600 1612.640 ;
        RECT 4.000 1609.240 2498.195 1611.240 ;
        RECT 4.400 1607.840 2495.600 1609.240 ;
        RECT 4.000 1605.840 2498.195 1607.840 ;
        RECT 4.400 1604.440 2495.600 1605.840 ;
        RECT 4.000 1602.440 2498.195 1604.440 ;
        RECT 4.400 1601.040 2495.600 1602.440 ;
        RECT 4.000 1599.040 2498.195 1601.040 ;
        RECT 4.400 1597.640 2495.600 1599.040 ;
        RECT 4.000 1595.640 2498.195 1597.640 ;
        RECT 4.400 1594.240 2495.600 1595.640 ;
        RECT 4.000 1592.240 2498.195 1594.240 ;
        RECT 4.400 1590.840 2495.600 1592.240 ;
        RECT 4.000 1588.840 2498.195 1590.840 ;
        RECT 4.400 1587.440 2495.600 1588.840 ;
        RECT 4.000 1585.440 2498.195 1587.440 ;
        RECT 4.400 1584.040 2495.600 1585.440 ;
        RECT 4.000 1582.040 2498.195 1584.040 ;
        RECT 4.400 1580.640 2498.195 1582.040 ;
        RECT 4.000 1578.640 2498.195 1580.640 ;
        RECT 4.400 1577.240 2495.600 1578.640 ;
        RECT 4.000 1575.240 2498.195 1577.240 ;
        RECT 4.400 1573.840 2495.600 1575.240 ;
        RECT 4.000 1571.840 2498.195 1573.840 ;
        RECT 4.400 1570.440 2495.600 1571.840 ;
        RECT 4.000 1568.440 2498.195 1570.440 ;
        RECT 4.000 1567.040 2495.600 1568.440 ;
        RECT 4.000 1565.040 2498.195 1567.040 ;
        RECT 4.400 1563.640 2495.600 1565.040 ;
        RECT 4.000 1561.640 2498.195 1563.640 ;
        RECT 4.400 1560.240 2495.600 1561.640 ;
        RECT 4.000 1558.240 2498.195 1560.240 ;
        RECT 4.400 1556.840 2495.600 1558.240 ;
        RECT 4.000 1554.840 2498.195 1556.840 ;
        RECT 4.400 1553.440 2495.600 1554.840 ;
        RECT 4.000 1551.440 2498.195 1553.440 ;
        RECT 4.400 1550.040 2495.600 1551.440 ;
        RECT 4.000 1548.040 2498.195 1550.040 ;
        RECT 4.400 1546.640 2495.600 1548.040 ;
        RECT 4.000 1544.640 2498.195 1546.640 ;
        RECT 4.400 1543.240 2495.600 1544.640 ;
        RECT 4.000 1541.240 2498.195 1543.240 ;
        RECT 4.400 1539.840 2495.600 1541.240 ;
        RECT 4.000 1537.840 2498.195 1539.840 ;
        RECT 4.400 1536.440 2495.600 1537.840 ;
        RECT 4.000 1534.440 2498.195 1536.440 ;
        RECT 4.400 1533.040 2495.600 1534.440 ;
        RECT 4.000 1531.040 2498.195 1533.040 ;
        RECT 4.400 1529.640 2495.600 1531.040 ;
        RECT 4.000 1527.640 2498.195 1529.640 ;
        RECT 4.400 1526.240 2498.195 1527.640 ;
        RECT 4.000 1524.240 2498.195 1526.240 ;
        RECT 4.400 1522.840 2495.600 1524.240 ;
        RECT 4.000 1520.840 2498.195 1522.840 ;
        RECT 4.400 1519.440 2495.600 1520.840 ;
        RECT 4.000 1517.440 2498.195 1519.440 ;
        RECT 4.400 1516.040 2495.600 1517.440 ;
        RECT 4.000 1514.040 2498.195 1516.040 ;
        RECT 4.000 1512.640 2495.600 1514.040 ;
        RECT 4.000 1510.640 2498.195 1512.640 ;
        RECT 4.400 1509.240 2495.600 1510.640 ;
        RECT 4.000 1507.240 2498.195 1509.240 ;
        RECT 4.400 1505.840 2495.600 1507.240 ;
        RECT 4.000 1503.840 2498.195 1505.840 ;
        RECT 4.400 1502.440 2495.600 1503.840 ;
        RECT 4.000 1500.440 2498.195 1502.440 ;
        RECT 4.400 1499.040 2495.600 1500.440 ;
        RECT 4.000 1497.040 2498.195 1499.040 ;
        RECT 4.400 1495.640 2495.600 1497.040 ;
        RECT 4.000 1493.640 2498.195 1495.640 ;
        RECT 4.400 1492.240 2495.600 1493.640 ;
        RECT 4.000 1490.240 2498.195 1492.240 ;
        RECT 4.400 1488.840 2495.600 1490.240 ;
        RECT 4.000 1486.840 2498.195 1488.840 ;
        RECT 4.400 1485.440 2495.600 1486.840 ;
        RECT 4.000 1483.440 2498.195 1485.440 ;
        RECT 4.400 1482.040 2495.600 1483.440 ;
        RECT 4.000 1480.040 2498.195 1482.040 ;
        RECT 4.400 1478.640 2495.600 1480.040 ;
        RECT 4.000 1476.640 2498.195 1478.640 ;
        RECT 4.400 1475.240 2495.600 1476.640 ;
        RECT 4.000 1473.240 2498.195 1475.240 ;
        RECT 4.400 1471.840 2498.195 1473.240 ;
        RECT 4.000 1469.840 2498.195 1471.840 ;
        RECT 4.400 1468.440 2495.600 1469.840 ;
        RECT 4.000 1466.440 2498.195 1468.440 ;
        RECT 4.400 1465.040 2495.600 1466.440 ;
        RECT 4.000 1463.040 2498.195 1465.040 ;
        RECT 4.000 1461.640 2495.600 1463.040 ;
        RECT 4.000 1459.640 2498.195 1461.640 ;
        RECT 4.400 1458.240 2495.600 1459.640 ;
        RECT 4.000 1456.240 2498.195 1458.240 ;
        RECT 4.400 1454.840 2495.600 1456.240 ;
        RECT 4.000 1452.840 2498.195 1454.840 ;
        RECT 4.400 1451.440 2495.600 1452.840 ;
        RECT 4.000 1449.440 2498.195 1451.440 ;
        RECT 4.400 1448.040 2495.600 1449.440 ;
        RECT 4.000 1446.040 2498.195 1448.040 ;
        RECT 4.400 1444.640 2495.600 1446.040 ;
        RECT 4.000 1442.640 2498.195 1444.640 ;
        RECT 4.400 1441.240 2495.600 1442.640 ;
        RECT 4.000 1439.240 2498.195 1441.240 ;
        RECT 4.400 1437.840 2495.600 1439.240 ;
        RECT 4.000 1435.840 2498.195 1437.840 ;
        RECT 4.400 1434.440 2495.600 1435.840 ;
        RECT 4.000 1432.440 2498.195 1434.440 ;
        RECT 4.400 1431.040 2495.600 1432.440 ;
        RECT 4.000 1429.040 2498.195 1431.040 ;
        RECT 4.400 1427.640 2495.600 1429.040 ;
        RECT 4.000 1425.640 2498.195 1427.640 ;
        RECT 4.400 1424.240 2495.600 1425.640 ;
        RECT 4.000 1422.240 2498.195 1424.240 ;
        RECT 4.400 1420.840 2495.600 1422.240 ;
        RECT 4.000 1418.840 2498.195 1420.840 ;
        RECT 4.400 1417.440 2498.195 1418.840 ;
        RECT 4.000 1415.440 2498.195 1417.440 ;
        RECT 4.400 1414.040 2495.600 1415.440 ;
        RECT 4.000 1412.040 2498.195 1414.040 ;
        RECT 4.400 1410.640 2495.600 1412.040 ;
        RECT 4.000 1408.640 2498.195 1410.640 ;
        RECT 4.000 1407.240 2495.600 1408.640 ;
        RECT 4.000 1405.240 2498.195 1407.240 ;
        RECT 4.400 1403.840 2495.600 1405.240 ;
        RECT 4.000 1401.840 2498.195 1403.840 ;
        RECT 4.400 1400.440 2495.600 1401.840 ;
        RECT 4.000 1398.440 2498.195 1400.440 ;
        RECT 4.400 1397.040 2495.600 1398.440 ;
        RECT 4.000 1395.040 2498.195 1397.040 ;
        RECT 4.400 1393.640 2495.600 1395.040 ;
        RECT 4.000 1391.640 2498.195 1393.640 ;
        RECT 4.400 1390.240 2495.600 1391.640 ;
        RECT 4.000 1388.240 2498.195 1390.240 ;
        RECT 4.400 1386.840 2495.600 1388.240 ;
        RECT 4.000 1384.840 2498.195 1386.840 ;
        RECT 4.400 1383.440 2495.600 1384.840 ;
        RECT 4.000 1381.440 2498.195 1383.440 ;
        RECT 4.400 1380.040 2495.600 1381.440 ;
        RECT 4.000 1378.040 2498.195 1380.040 ;
        RECT 4.400 1376.640 2495.600 1378.040 ;
        RECT 4.000 1374.640 2498.195 1376.640 ;
        RECT 4.400 1373.240 2495.600 1374.640 ;
        RECT 4.000 1371.240 2498.195 1373.240 ;
        RECT 4.400 1369.840 2495.600 1371.240 ;
        RECT 4.000 1367.840 2498.195 1369.840 ;
        RECT 4.400 1366.440 2495.600 1367.840 ;
        RECT 4.000 1364.440 2498.195 1366.440 ;
        RECT 4.400 1363.040 2498.195 1364.440 ;
        RECT 4.000 1361.040 2498.195 1363.040 ;
        RECT 4.400 1359.640 2495.600 1361.040 ;
        RECT 4.000 1357.640 2498.195 1359.640 ;
        RECT 4.400 1356.240 2495.600 1357.640 ;
        RECT 4.000 1354.240 2498.195 1356.240 ;
        RECT 4.000 1352.840 2495.600 1354.240 ;
        RECT 4.000 1350.840 2498.195 1352.840 ;
        RECT 4.400 1349.440 2495.600 1350.840 ;
        RECT 4.000 1347.440 2498.195 1349.440 ;
        RECT 4.400 1346.040 2495.600 1347.440 ;
        RECT 4.000 1344.040 2498.195 1346.040 ;
        RECT 4.400 1342.640 2495.600 1344.040 ;
        RECT 4.000 1340.640 2498.195 1342.640 ;
        RECT 4.400 1339.240 2495.600 1340.640 ;
        RECT 4.000 1337.240 2498.195 1339.240 ;
        RECT 4.400 1335.840 2495.600 1337.240 ;
        RECT 4.000 1333.840 2498.195 1335.840 ;
        RECT 4.400 1332.440 2495.600 1333.840 ;
        RECT 4.000 1330.440 2498.195 1332.440 ;
        RECT 4.400 1329.040 2495.600 1330.440 ;
        RECT 4.000 1327.040 2498.195 1329.040 ;
        RECT 4.400 1325.640 2495.600 1327.040 ;
        RECT 4.000 1323.640 2498.195 1325.640 ;
        RECT 4.400 1322.240 2495.600 1323.640 ;
        RECT 4.000 1320.240 2498.195 1322.240 ;
        RECT 4.400 1318.840 2495.600 1320.240 ;
        RECT 4.000 1316.840 2498.195 1318.840 ;
        RECT 4.400 1315.440 2495.600 1316.840 ;
        RECT 4.000 1313.440 2498.195 1315.440 ;
        RECT 4.400 1312.040 2495.600 1313.440 ;
        RECT 4.000 1310.040 2498.195 1312.040 ;
        RECT 4.400 1308.640 2498.195 1310.040 ;
        RECT 4.000 1306.640 2498.195 1308.640 ;
        RECT 4.400 1305.240 2495.600 1306.640 ;
        RECT 4.000 1303.240 2498.195 1305.240 ;
        RECT 4.400 1301.840 2495.600 1303.240 ;
        RECT 4.000 1299.840 2498.195 1301.840 ;
        RECT 4.000 1298.440 2495.600 1299.840 ;
        RECT 4.000 1296.440 2498.195 1298.440 ;
        RECT 4.400 1295.040 2495.600 1296.440 ;
        RECT 4.000 1293.040 2498.195 1295.040 ;
        RECT 4.400 1291.640 2495.600 1293.040 ;
        RECT 4.000 1289.640 2498.195 1291.640 ;
        RECT 4.400 1288.240 2495.600 1289.640 ;
        RECT 4.000 1286.240 2498.195 1288.240 ;
        RECT 4.400 1284.840 2495.600 1286.240 ;
        RECT 4.000 1282.840 2498.195 1284.840 ;
        RECT 4.400 1281.440 2495.600 1282.840 ;
        RECT 4.000 1279.440 2498.195 1281.440 ;
        RECT 4.400 1278.040 2495.600 1279.440 ;
        RECT 4.000 1276.040 2498.195 1278.040 ;
        RECT 4.400 1274.640 2495.600 1276.040 ;
        RECT 4.000 1272.640 2498.195 1274.640 ;
        RECT 4.400 1271.240 2495.600 1272.640 ;
        RECT 4.000 1269.240 2498.195 1271.240 ;
        RECT 4.400 1267.840 2495.600 1269.240 ;
        RECT 4.000 1265.840 2498.195 1267.840 ;
        RECT 4.400 1264.440 2495.600 1265.840 ;
        RECT 4.000 1262.440 2498.195 1264.440 ;
        RECT 4.400 1261.040 2495.600 1262.440 ;
        RECT 4.000 1259.040 2498.195 1261.040 ;
        RECT 4.400 1257.640 2495.600 1259.040 ;
        RECT 4.000 1255.640 2498.195 1257.640 ;
        RECT 4.400 1254.240 2498.195 1255.640 ;
        RECT 4.000 1252.240 2498.195 1254.240 ;
        RECT 4.400 1250.840 2495.600 1252.240 ;
        RECT 4.000 1248.840 2498.195 1250.840 ;
        RECT 4.400 1247.440 2495.600 1248.840 ;
        RECT 4.000 1245.440 2498.195 1247.440 ;
        RECT 4.000 1244.040 2495.600 1245.440 ;
        RECT 4.000 1242.040 2498.195 1244.040 ;
        RECT 4.400 1240.640 2495.600 1242.040 ;
        RECT 4.000 1238.640 2498.195 1240.640 ;
        RECT 4.400 1237.240 2495.600 1238.640 ;
        RECT 4.000 1235.240 2498.195 1237.240 ;
        RECT 4.400 1233.840 2495.600 1235.240 ;
        RECT 4.000 1231.840 2498.195 1233.840 ;
        RECT 4.400 1230.440 2495.600 1231.840 ;
        RECT 4.000 1228.440 2498.195 1230.440 ;
        RECT 4.400 1227.040 2495.600 1228.440 ;
        RECT 4.000 1225.040 2498.195 1227.040 ;
        RECT 4.400 1223.640 2495.600 1225.040 ;
        RECT 4.000 1221.640 2498.195 1223.640 ;
        RECT 4.400 1220.240 2495.600 1221.640 ;
        RECT 4.000 1218.240 2498.195 1220.240 ;
        RECT 4.400 1216.840 2495.600 1218.240 ;
        RECT 4.000 1214.840 2498.195 1216.840 ;
        RECT 4.400 1213.440 2495.600 1214.840 ;
        RECT 4.000 1211.440 2498.195 1213.440 ;
        RECT 4.400 1210.040 2495.600 1211.440 ;
        RECT 4.000 1208.040 2498.195 1210.040 ;
        RECT 4.400 1206.640 2495.600 1208.040 ;
        RECT 4.000 1204.640 2498.195 1206.640 ;
        RECT 4.400 1203.240 2495.600 1204.640 ;
        RECT 4.000 1201.240 2498.195 1203.240 ;
        RECT 4.400 1199.840 2498.195 1201.240 ;
        RECT 4.000 1197.840 2498.195 1199.840 ;
        RECT 4.400 1196.440 2495.600 1197.840 ;
        RECT 4.000 1194.440 2498.195 1196.440 ;
        RECT 4.400 1193.040 2495.600 1194.440 ;
        RECT 4.000 1191.040 2498.195 1193.040 ;
        RECT 4.000 1189.640 2495.600 1191.040 ;
        RECT 4.000 1187.640 2498.195 1189.640 ;
        RECT 4.400 1186.240 2495.600 1187.640 ;
        RECT 4.000 1184.240 2498.195 1186.240 ;
        RECT 4.400 1182.840 2495.600 1184.240 ;
        RECT 4.000 1180.840 2498.195 1182.840 ;
        RECT 4.400 1179.440 2495.600 1180.840 ;
        RECT 4.000 1177.440 2498.195 1179.440 ;
        RECT 4.400 1176.040 2495.600 1177.440 ;
        RECT 4.000 1174.040 2498.195 1176.040 ;
        RECT 4.400 1172.640 2495.600 1174.040 ;
        RECT 4.000 1170.640 2498.195 1172.640 ;
        RECT 4.400 1169.240 2495.600 1170.640 ;
        RECT 4.000 1167.240 2498.195 1169.240 ;
        RECT 4.400 1165.840 2495.600 1167.240 ;
        RECT 4.000 1163.840 2498.195 1165.840 ;
        RECT 4.400 1162.440 2495.600 1163.840 ;
        RECT 4.000 1160.440 2498.195 1162.440 ;
        RECT 4.400 1159.040 2495.600 1160.440 ;
        RECT 4.000 1157.040 2498.195 1159.040 ;
        RECT 4.400 1155.640 2495.600 1157.040 ;
        RECT 4.000 1153.640 2498.195 1155.640 ;
        RECT 4.400 1152.240 2495.600 1153.640 ;
        RECT 4.000 1150.240 2498.195 1152.240 ;
        RECT 4.400 1148.840 2495.600 1150.240 ;
        RECT 4.000 1146.840 2498.195 1148.840 ;
        RECT 4.400 1145.440 2498.195 1146.840 ;
        RECT 4.000 1143.440 2498.195 1145.440 ;
        RECT 4.400 1142.040 2495.600 1143.440 ;
        RECT 4.000 1140.040 2498.195 1142.040 ;
        RECT 4.400 1138.640 2495.600 1140.040 ;
        RECT 4.000 1136.640 2498.195 1138.640 ;
        RECT 4.000 1135.240 2495.600 1136.640 ;
        RECT 4.000 1133.240 2498.195 1135.240 ;
        RECT 4.400 1131.840 2495.600 1133.240 ;
        RECT 4.000 1129.840 2498.195 1131.840 ;
        RECT 4.400 1128.440 2495.600 1129.840 ;
        RECT 4.000 1126.440 2498.195 1128.440 ;
        RECT 4.400 1125.040 2495.600 1126.440 ;
        RECT 4.000 1123.040 2498.195 1125.040 ;
        RECT 4.400 1121.640 2495.600 1123.040 ;
        RECT 4.000 1119.640 2498.195 1121.640 ;
        RECT 4.400 1118.240 2495.600 1119.640 ;
        RECT 4.000 1116.240 2498.195 1118.240 ;
        RECT 4.400 1114.840 2495.600 1116.240 ;
        RECT 4.000 1112.840 2498.195 1114.840 ;
        RECT 4.400 1111.440 2495.600 1112.840 ;
        RECT 4.000 1109.440 2498.195 1111.440 ;
        RECT 4.400 1108.040 2495.600 1109.440 ;
        RECT 4.000 1106.040 2498.195 1108.040 ;
        RECT 4.400 1104.640 2495.600 1106.040 ;
        RECT 4.000 1102.640 2498.195 1104.640 ;
        RECT 4.400 1101.240 2495.600 1102.640 ;
        RECT 4.000 1099.240 2498.195 1101.240 ;
        RECT 4.400 1097.840 2495.600 1099.240 ;
        RECT 4.000 1095.840 2498.195 1097.840 ;
        RECT 4.400 1094.440 2495.600 1095.840 ;
        RECT 4.000 1092.440 2498.195 1094.440 ;
        RECT 4.400 1091.040 2498.195 1092.440 ;
        RECT 4.000 1089.040 2498.195 1091.040 ;
        RECT 4.400 1087.640 2495.600 1089.040 ;
        RECT 4.000 1085.640 2498.195 1087.640 ;
        RECT 4.400 1084.240 2495.600 1085.640 ;
        RECT 4.000 1082.240 2498.195 1084.240 ;
        RECT 4.000 1080.840 2495.600 1082.240 ;
        RECT 4.000 1078.840 2498.195 1080.840 ;
        RECT 4.400 1077.440 2495.600 1078.840 ;
        RECT 4.000 1075.440 2498.195 1077.440 ;
        RECT 4.400 1074.040 2495.600 1075.440 ;
        RECT 4.000 1072.040 2498.195 1074.040 ;
        RECT 4.400 1070.640 2495.600 1072.040 ;
        RECT 4.000 1068.640 2498.195 1070.640 ;
        RECT 4.400 1067.240 2495.600 1068.640 ;
        RECT 4.000 1065.240 2498.195 1067.240 ;
        RECT 4.400 1063.840 2495.600 1065.240 ;
        RECT 4.000 1061.840 2498.195 1063.840 ;
        RECT 4.400 1060.440 2495.600 1061.840 ;
        RECT 4.000 1058.440 2498.195 1060.440 ;
        RECT 4.400 1057.040 2495.600 1058.440 ;
        RECT 4.000 1055.040 2498.195 1057.040 ;
        RECT 4.400 1053.640 2495.600 1055.040 ;
        RECT 4.000 1051.640 2498.195 1053.640 ;
        RECT 4.400 1050.240 2495.600 1051.640 ;
        RECT 4.000 1048.240 2498.195 1050.240 ;
        RECT 4.400 1046.840 2495.600 1048.240 ;
        RECT 4.000 1044.840 2498.195 1046.840 ;
        RECT 4.400 1043.440 2495.600 1044.840 ;
        RECT 4.000 1041.440 2498.195 1043.440 ;
        RECT 4.400 1040.040 2495.600 1041.440 ;
        RECT 4.000 1038.040 2498.195 1040.040 ;
        RECT 4.400 1036.640 2498.195 1038.040 ;
        RECT 4.000 1034.640 2498.195 1036.640 ;
        RECT 4.400 1033.240 2495.600 1034.640 ;
        RECT 4.000 1031.240 2498.195 1033.240 ;
        RECT 4.400 1029.840 2495.600 1031.240 ;
        RECT 4.000 1027.840 2498.195 1029.840 ;
        RECT 4.000 1026.440 2495.600 1027.840 ;
        RECT 4.000 1024.440 2498.195 1026.440 ;
        RECT 4.400 1023.040 2495.600 1024.440 ;
        RECT 4.000 1021.040 2498.195 1023.040 ;
        RECT 4.400 1019.640 2495.600 1021.040 ;
        RECT 4.000 1017.640 2498.195 1019.640 ;
        RECT 4.400 1016.240 2495.600 1017.640 ;
        RECT 4.000 1014.240 2498.195 1016.240 ;
        RECT 4.400 1012.840 2495.600 1014.240 ;
        RECT 4.000 1010.840 2498.195 1012.840 ;
        RECT 4.400 1009.440 2495.600 1010.840 ;
        RECT 4.000 1007.440 2498.195 1009.440 ;
        RECT 4.400 1006.040 2495.600 1007.440 ;
        RECT 4.000 1004.040 2498.195 1006.040 ;
        RECT 4.400 1002.640 2495.600 1004.040 ;
        RECT 4.000 1000.640 2498.195 1002.640 ;
        RECT 4.400 999.240 2495.600 1000.640 ;
        RECT 4.000 997.240 2498.195 999.240 ;
        RECT 4.400 995.840 2495.600 997.240 ;
        RECT 4.000 993.840 2498.195 995.840 ;
        RECT 4.400 992.440 2495.600 993.840 ;
        RECT 4.000 990.440 2498.195 992.440 ;
        RECT 4.400 989.040 2495.600 990.440 ;
        RECT 4.000 987.040 2498.195 989.040 ;
        RECT 4.400 985.640 2498.195 987.040 ;
        RECT 4.000 983.640 2498.195 985.640 ;
        RECT 4.400 982.240 2495.600 983.640 ;
        RECT 4.000 980.240 2498.195 982.240 ;
        RECT 4.400 978.840 2495.600 980.240 ;
        RECT 4.000 976.840 2498.195 978.840 ;
        RECT 4.400 975.440 2495.600 976.840 ;
        RECT 4.000 973.440 2498.195 975.440 ;
        RECT 4.000 972.040 2495.600 973.440 ;
        RECT 4.000 970.040 2498.195 972.040 ;
        RECT 4.400 968.640 2495.600 970.040 ;
        RECT 4.000 966.640 2498.195 968.640 ;
        RECT 4.400 965.240 2495.600 966.640 ;
        RECT 4.000 963.240 2498.195 965.240 ;
        RECT 4.400 961.840 2495.600 963.240 ;
        RECT 4.000 959.840 2498.195 961.840 ;
        RECT 4.400 958.440 2495.600 959.840 ;
        RECT 4.000 956.440 2498.195 958.440 ;
        RECT 4.400 955.040 2495.600 956.440 ;
        RECT 4.000 953.040 2498.195 955.040 ;
        RECT 4.400 951.640 2495.600 953.040 ;
        RECT 4.000 949.640 2498.195 951.640 ;
        RECT 4.400 948.240 2495.600 949.640 ;
        RECT 4.000 946.240 2498.195 948.240 ;
        RECT 4.400 944.840 2495.600 946.240 ;
        RECT 4.000 942.840 2498.195 944.840 ;
        RECT 4.400 941.440 2495.600 942.840 ;
        RECT 4.000 939.440 2498.195 941.440 ;
        RECT 4.400 938.040 2495.600 939.440 ;
        RECT 4.000 936.040 2498.195 938.040 ;
        RECT 4.400 934.640 2495.600 936.040 ;
        RECT 4.000 932.640 2498.195 934.640 ;
        RECT 4.400 931.240 2498.195 932.640 ;
        RECT 4.000 929.240 2498.195 931.240 ;
        RECT 4.400 927.840 2495.600 929.240 ;
        RECT 4.000 925.840 2498.195 927.840 ;
        RECT 4.400 924.440 2495.600 925.840 ;
        RECT 4.000 922.440 2498.195 924.440 ;
        RECT 4.400 921.040 2495.600 922.440 ;
        RECT 4.000 919.040 2498.195 921.040 ;
        RECT 4.000 917.640 2495.600 919.040 ;
        RECT 4.000 915.640 2498.195 917.640 ;
        RECT 4.400 914.240 2495.600 915.640 ;
        RECT 4.000 912.240 2498.195 914.240 ;
        RECT 4.400 910.840 2495.600 912.240 ;
        RECT 4.000 908.840 2498.195 910.840 ;
        RECT 4.400 907.440 2495.600 908.840 ;
        RECT 4.000 905.440 2498.195 907.440 ;
        RECT 4.400 904.040 2495.600 905.440 ;
        RECT 4.000 902.040 2498.195 904.040 ;
        RECT 4.400 900.640 2495.600 902.040 ;
        RECT 4.000 898.640 2498.195 900.640 ;
        RECT 4.400 897.240 2495.600 898.640 ;
        RECT 4.000 895.240 2498.195 897.240 ;
        RECT 4.400 893.840 2495.600 895.240 ;
        RECT 4.000 891.840 2498.195 893.840 ;
        RECT 4.400 890.440 2495.600 891.840 ;
        RECT 4.000 888.440 2498.195 890.440 ;
        RECT 4.400 887.040 2495.600 888.440 ;
        RECT 4.000 885.040 2498.195 887.040 ;
        RECT 4.400 883.640 2495.600 885.040 ;
        RECT 4.000 881.640 2498.195 883.640 ;
        RECT 4.400 880.240 2495.600 881.640 ;
        RECT 4.000 878.240 2498.195 880.240 ;
        RECT 4.400 876.840 2498.195 878.240 ;
        RECT 4.000 874.840 2498.195 876.840 ;
        RECT 4.400 873.440 2495.600 874.840 ;
        RECT 4.000 871.440 2498.195 873.440 ;
        RECT 4.400 870.040 2495.600 871.440 ;
        RECT 4.000 868.040 2498.195 870.040 ;
        RECT 4.400 866.640 2495.600 868.040 ;
        RECT 4.000 864.640 2498.195 866.640 ;
        RECT 4.000 863.240 2495.600 864.640 ;
        RECT 4.000 861.240 2498.195 863.240 ;
        RECT 4.400 859.840 2495.600 861.240 ;
        RECT 4.000 857.840 2498.195 859.840 ;
        RECT 4.400 856.440 2495.600 857.840 ;
        RECT 4.000 854.440 2498.195 856.440 ;
        RECT 4.400 853.040 2495.600 854.440 ;
        RECT 4.000 851.040 2498.195 853.040 ;
        RECT 4.400 849.640 2495.600 851.040 ;
        RECT 4.000 847.640 2498.195 849.640 ;
        RECT 4.400 846.240 2495.600 847.640 ;
        RECT 4.000 844.240 2498.195 846.240 ;
        RECT 4.400 842.840 2495.600 844.240 ;
        RECT 4.000 840.840 2498.195 842.840 ;
        RECT 4.400 839.440 2495.600 840.840 ;
        RECT 4.000 837.440 2498.195 839.440 ;
        RECT 4.400 836.040 2495.600 837.440 ;
        RECT 4.000 834.040 2498.195 836.040 ;
        RECT 4.400 832.640 2495.600 834.040 ;
        RECT 4.000 830.640 2498.195 832.640 ;
        RECT 4.400 829.240 2495.600 830.640 ;
        RECT 4.000 827.240 2498.195 829.240 ;
        RECT 4.400 825.840 2495.600 827.240 ;
        RECT 4.000 823.840 2498.195 825.840 ;
        RECT 4.400 822.440 2498.195 823.840 ;
        RECT 4.000 820.440 2498.195 822.440 ;
        RECT 4.400 819.040 2495.600 820.440 ;
        RECT 4.000 817.040 2498.195 819.040 ;
        RECT 4.400 815.640 2495.600 817.040 ;
        RECT 4.000 813.640 2498.195 815.640 ;
        RECT 4.400 812.240 2495.600 813.640 ;
        RECT 4.000 810.240 2498.195 812.240 ;
        RECT 4.000 808.840 2495.600 810.240 ;
        RECT 4.000 806.840 2498.195 808.840 ;
        RECT 4.400 805.440 2495.600 806.840 ;
        RECT 4.000 803.440 2498.195 805.440 ;
        RECT 4.400 802.040 2495.600 803.440 ;
        RECT 4.000 800.040 2498.195 802.040 ;
        RECT 4.400 798.640 2495.600 800.040 ;
        RECT 4.000 796.640 2498.195 798.640 ;
        RECT 4.400 795.240 2495.600 796.640 ;
        RECT 4.000 793.240 2498.195 795.240 ;
        RECT 4.400 791.840 2495.600 793.240 ;
        RECT 4.000 789.840 2498.195 791.840 ;
        RECT 4.400 788.440 2495.600 789.840 ;
        RECT 4.000 786.440 2498.195 788.440 ;
        RECT 4.400 785.040 2495.600 786.440 ;
        RECT 4.000 783.040 2498.195 785.040 ;
        RECT 4.400 781.640 2495.600 783.040 ;
        RECT 4.000 779.640 2498.195 781.640 ;
        RECT 4.400 778.240 2495.600 779.640 ;
        RECT 4.000 776.240 2498.195 778.240 ;
        RECT 4.400 774.840 2495.600 776.240 ;
        RECT 4.000 772.840 2498.195 774.840 ;
        RECT 4.400 771.440 2495.600 772.840 ;
        RECT 4.000 769.440 2498.195 771.440 ;
        RECT 4.400 768.040 2498.195 769.440 ;
        RECT 4.000 766.040 2498.195 768.040 ;
        RECT 4.400 764.640 2495.600 766.040 ;
        RECT 4.000 762.640 2498.195 764.640 ;
        RECT 4.400 761.240 2495.600 762.640 ;
        RECT 4.000 759.240 2498.195 761.240 ;
        RECT 4.400 757.840 2495.600 759.240 ;
        RECT 4.000 755.840 2498.195 757.840 ;
        RECT 4.000 754.440 2495.600 755.840 ;
        RECT 4.000 752.440 2498.195 754.440 ;
        RECT 4.400 751.040 2495.600 752.440 ;
        RECT 4.000 749.040 2498.195 751.040 ;
        RECT 4.400 747.640 2495.600 749.040 ;
        RECT 4.000 745.640 2498.195 747.640 ;
        RECT 4.400 744.240 2495.600 745.640 ;
        RECT 4.000 742.240 2498.195 744.240 ;
        RECT 4.400 740.840 2495.600 742.240 ;
        RECT 4.000 738.840 2498.195 740.840 ;
        RECT 4.400 737.440 2495.600 738.840 ;
        RECT 4.000 735.440 2498.195 737.440 ;
        RECT 4.400 734.040 2495.600 735.440 ;
        RECT 4.000 732.040 2498.195 734.040 ;
        RECT 4.400 730.640 2495.600 732.040 ;
        RECT 4.000 728.640 2498.195 730.640 ;
        RECT 4.400 727.240 2495.600 728.640 ;
        RECT 4.000 725.240 2498.195 727.240 ;
        RECT 4.400 723.840 2495.600 725.240 ;
        RECT 4.000 721.840 2498.195 723.840 ;
        RECT 4.400 720.440 2495.600 721.840 ;
        RECT 4.000 718.440 2498.195 720.440 ;
        RECT 4.400 717.040 2495.600 718.440 ;
        RECT 4.000 715.040 2498.195 717.040 ;
        RECT 4.400 713.640 2498.195 715.040 ;
        RECT 4.000 711.640 2498.195 713.640 ;
        RECT 4.400 710.240 2495.600 711.640 ;
        RECT 4.000 708.240 2498.195 710.240 ;
        RECT 4.400 706.840 2495.600 708.240 ;
        RECT 4.000 704.840 2498.195 706.840 ;
        RECT 4.000 703.440 2495.600 704.840 ;
        RECT 4.000 701.440 2498.195 703.440 ;
        RECT 4.400 700.040 2495.600 701.440 ;
        RECT 4.000 698.040 2498.195 700.040 ;
        RECT 4.400 696.640 2495.600 698.040 ;
        RECT 4.000 694.640 2498.195 696.640 ;
        RECT 4.400 693.240 2495.600 694.640 ;
        RECT 4.000 691.240 2498.195 693.240 ;
        RECT 4.400 689.840 2495.600 691.240 ;
        RECT 4.000 687.840 2498.195 689.840 ;
        RECT 4.400 686.440 2495.600 687.840 ;
        RECT 4.000 684.440 2498.195 686.440 ;
        RECT 4.400 683.040 2495.600 684.440 ;
        RECT 4.000 681.040 2498.195 683.040 ;
        RECT 4.400 679.640 2495.600 681.040 ;
        RECT 4.000 677.640 2498.195 679.640 ;
        RECT 4.400 676.240 2495.600 677.640 ;
        RECT 4.000 674.240 2498.195 676.240 ;
        RECT 4.400 672.840 2495.600 674.240 ;
        RECT 4.000 670.840 2498.195 672.840 ;
        RECT 4.400 669.440 2495.600 670.840 ;
        RECT 4.000 667.440 2498.195 669.440 ;
        RECT 4.400 666.040 2495.600 667.440 ;
        RECT 4.000 664.040 2498.195 666.040 ;
        RECT 4.400 662.640 2495.600 664.040 ;
        RECT 4.000 660.640 2498.195 662.640 ;
        RECT 4.400 659.240 2498.195 660.640 ;
        RECT 4.000 657.240 2498.195 659.240 ;
        RECT 4.400 655.840 2495.600 657.240 ;
        RECT 4.000 653.840 2498.195 655.840 ;
        RECT 4.400 652.440 2495.600 653.840 ;
        RECT 4.000 650.440 2498.195 652.440 ;
        RECT 4.000 649.040 2495.600 650.440 ;
        RECT 4.000 647.040 2498.195 649.040 ;
        RECT 4.400 645.640 2495.600 647.040 ;
        RECT 4.000 643.640 2498.195 645.640 ;
        RECT 4.400 642.240 2495.600 643.640 ;
        RECT 4.000 640.240 2498.195 642.240 ;
        RECT 4.400 638.840 2495.600 640.240 ;
        RECT 4.000 636.840 2498.195 638.840 ;
        RECT 4.400 635.440 2495.600 636.840 ;
        RECT 4.000 633.440 2498.195 635.440 ;
        RECT 4.400 632.040 2495.600 633.440 ;
        RECT 4.000 630.040 2498.195 632.040 ;
        RECT 4.400 628.640 2495.600 630.040 ;
        RECT 4.000 626.640 2498.195 628.640 ;
        RECT 4.400 625.240 2495.600 626.640 ;
        RECT 4.000 623.240 2498.195 625.240 ;
        RECT 4.400 621.840 2495.600 623.240 ;
        RECT 4.000 619.840 2498.195 621.840 ;
        RECT 4.400 618.440 2495.600 619.840 ;
        RECT 4.000 616.440 2498.195 618.440 ;
        RECT 4.400 615.040 2495.600 616.440 ;
        RECT 4.000 613.040 2498.195 615.040 ;
        RECT 4.400 611.640 2495.600 613.040 ;
        RECT 4.000 609.640 2498.195 611.640 ;
        RECT 4.400 608.240 2495.600 609.640 ;
        RECT 4.000 606.240 2498.195 608.240 ;
        RECT 4.400 604.840 2498.195 606.240 ;
        RECT 4.000 602.840 2498.195 604.840 ;
        RECT 4.400 601.440 2495.600 602.840 ;
        RECT 4.000 599.440 2498.195 601.440 ;
        RECT 4.400 598.040 2495.600 599.440 ;
        RECT 4.000 596.040 2498.195 598.040 ;
        RECT 4.000 594.640 2495.600 596.040 ;
        RECT 4.000 592.640 2498.195 594.640 ;
        RECT 4.400 591.240 2495.600 592.640 ;
        RECT 4.000 589.240 2498.195 591.240 ;
        RECT 4.400 587.840 2495.600 589.240 ;
        RECT 4.000 585.840 2498.195 587.840 ;
        RECT 4.400 584.440 2495.600 585.840 ;
        RECT 4.000 582.440 2498.195 584.440 ;
        RECT 4.400 581.040 2495.600 582.440 ;
        RECT 4.000 579.040 2498.195 581.040 ;
        RECT 4.400 577.640 2495.600 579.040 ;
        RECT 4.000 575.640 2498.195 577.640 ;
        RECT 4.400 574.240 2495.600 575.640 ;
        RECT 4.000 572.240 2498.195 574.240 ;
        RECT 4.400 570.840 2495.600 572.240 ;
        RECT 4.000 568.840 2498.195 570.840 ;
        RECT 4.400 567.440 2495.600 568.840 ;
        RECT 4.000 565.440 2498.195 567.440 ;
        RECT 4.400 564.040 2495.600 565.440 ;
        RECT 4.000 562.040 2498.195 564.040 ;
        RECT 4.400 560.640 2495.600 562.040 ;
        RECT 4.000 558.640 2498.195 560.640 ;
        RECT 4.400 557.240 2495.600 558.640 ;
        RECT 4.000 555.240 2498.195 557.240 ;
        RECT 4.400 553.840 2495.600 555.240 ;
        RECT 4.000 551.840 2498.195 553.840 ;
        RECT 4.400 550.440 2498.195 551.840 ;
        RECT 4.000 548.440 2498.195 550.440 ;
        RECT 4.400 547.040 2495.600 548.440 ;
        RECT 4.000 545.040 2498.195 547.040 ;
        RECT 4.400 543.640 2495.600 545.040 ;
        RECT 4.000 541.640 2498.195 543.640 ;
        RECT 4.000 540.240 2495.600 541.640 ;
        RECT 4.000 538.240 2498.195 540.240 ;
        RECT 4.400 536.840 2495.600 538.240 ;
        RECT 4.000 534.840 2498.195 536.840 ;
        RECT 4.400 533.440 2495.600 534.840 ;
        RECT 4.000 531.440 2498.195 533.440 ;
        RECT 4.400 530.040 2495.600 531.440 ;
        RECT 4.000 528.040 2498.195 530.040 ;
        RECT 4.400 526.640 2495.600 528.040 ;
        RECT 4.000 524.640 2498.195 526.640 ;
        RECT 4.400 523.240 2495.600 524.640 ;
        RECT 4.000 521.240 2498.195 523.240 ;
        RECT 4.400 519.840 2495.600 521.240 ;
        RECT 4.000 517.840 2498.195 519.840 ;
        RECT 4.400 516.440 2495.600 517.840 ;
        RECT 4.000 514.440 2498.195 516.440 ;
        RECT 4.400 513.040 2495.600 514.440 ;
        RECT 4.000 511.040 2498.195 513.040 ;
        RECT 4.400 509.640 2495.600 511.040 ;
        RECT 4.000 507.640 2498.195 509.640 ;
        RECT 4.400 506.240 2495.600 507.640 ;
        RECT 4.000 504.240 2498.195 506.240 ;
        RECT 4.400 502.840 2495.600 504.240 ;
        RECT 4.000 500.840 2498.195 502.840 ;
        RECT 4.400 499.440 2495.600 500.840 ;
        RECT 4.000 497.440 2498.195 499.440 ;
        RECT 4.400 496.040 2498.195 497.440 ;
        RECT 4.000 494.040 2498.195 496.040 ;
        RECT 4.400 492.640 2495.600 494.040 ;
        RECT 4.000 490.640 2498.195 492.640 ;
        RECT 4.400 489.240 2495.600 490.640 ;
        RECT 4.000 487.240 2498.195 489.240 ;
        RECT 4.000 485.840 2495.600 487.240 ;
        RECT 4.000 483.840 2498.195 485.840 ;
        RECT 4.400 482.440 2495.600 483.840 ;
        RECT 4.000 480.440 2498.195 482.440 ;
        RECT 4.400 479.040 2495.600 480.440 ;
        RECT 4.000 477.040 2498.195 479.040 ;
        RECT 4.400 475.640 2495.600 477.040 ;
        RECT 4.000 473.640 2498.195 475.640 ;
        RECT 4.400 472.240 2495.600 473.640 ;
        RECT 4.000 470.240 2498.195 472.240 ;
        RECT 4.400 468.840 2495.600 470.240 ;
        RECT 4.000 466.840 2498.195 468.840 ;
        RECT 4.400 465.440 2495.600 466.840 ;
        RECT 4.000 463.440 2498.195 465.440 ;
        RECT 4.400 462.040 2495.600 463.440 ;
        RECT 4.000 460.040 2498.195 462.040 ;
        RECT 4.400 458.640 2495.600 460.040 ;
        RECT 4.000 456.640 2498.195 458.640 ;
        RECT 4.400 455.240 2495.600 456.640 ;
        RECT 4.000 453.240 2498.195 455.240 ;
        RECT 4.400 451.840 2495.600 453.240 ;
        RECT 4.000 449.840 2498.195 451.840 ;
        RECT 4.400 448.440 2495.600 449.840 ;
        RECT 4.000 446.440 2498.195 448.440 ;
        RECT 4.400 445.040 2495.600 446.440 ;
        RECT 4.000 443.040 2498.195 445.040 ;
        RECT 4.400 441.640 2498.195 443.040 ;
        RECT 4.000 439.640 2498.195 441.640 ;
        RECT 4.400 438.240 2495.600 439.640 ;
        RECT 4.000 436.240 2498.195 438.240 ;
        RECT 4.400 434.840 2495.600 436.240 ;
        RECT 4.000 432.840 2498.195 434.840 ;
        RECT 4.000 431.440 2495.600 432.840 ;
        RECT 4.000 429.440 2498.195 431.440 ;
        RECT 4.400 428.040 2495.600 429.440 ;
        RECT 4.000 426.040 2498.195 428.040 ;
        RECT 4.400 424.640 2495.600 426.040 ;
        RECT 4.000 422.640 2498.195 424.640 ;
        RECT 4.400 421.240 2495.600 422.640 ;
        RECT 4.000 419.240 2498.195 421.240 ;
        RECT 4.400 417.840 2495.600 419.240 ;
        RECT 4.000 415.840 2498.195 417.840 ;
        RECT 4.400 414.440 2495.600 415.840 ;
        RECT 4.000 412.440 2498.195 414.440 ;
        RECT 4.400 411.040 2495.600 412.440 ;
        RECT 4.000 409.040 2498.195 411.040 ;
        RECT 4.400 407.640 2495.600 409.040 ;
        RECT 4.000 405.640 2498.195 407.640 ;
        RECT 4.400 404.240 2495.600 405.640 ;
        RECT 4.000 402.240 2498.195 404.240 ;
        RECT 4.400 400.840 2495.600 402.240 ;
        RECT 4.000 398.840 2498.195 400.840 ;
        RECT 4.400 397.440 2495.600 398.840 ;
        RECT 4.000 395.440 2498.195 397.440 ;
        RECT 4.400 394.040 2495.600 395.440 ;
        RECT 4.000 392.040 2498.195 394.040 ;
        RECT 4.400 390.640 2495.600 392.040 ;
        RECT 4.000 388.640 2498.195 390.640 ;
        RECT 4.400 387.240 2498.195 388.640 ;
        RECT 4.000 385.240 2498.195 387.240 ;
        RECT 4.400 383.840 2495.600 385.240 ;
        RECT 4.000 381.840 2498.195 383.840 ;
        RECT 4.400 380.440 2495.600 381.840 ;
        RECT 4.000 378.440 2498.195 380.440 ;
        RECT 4.000 377.040 2495.600 378.440 ;
        RECT 4.000 375.040 2498.195 377.040 ;
        RECT 4.400 373.640 2495.600 375.040 ;
        RECT 4.000 371.640 2498.195 373.640 ;
        RECT 4.400 370.240 2495.600 371.640 ;
        RECT 4.000 368.240 2498.195 370.240 ;
        RECT 4.400 366.840 2495.600 368.240 ;
        RECT 4.000 364.840 2498.195 366.840 ;
        RECT 4.400 363.440 2495.600 364.840 ;
        RECT 4.000 361.440 2498.195 363.440 ;
        RECT 4.400 360.040 2495.600 361.440 ;
        RECT 4.000 358.040 2498.195 360.040 ;
        RECT 4.400 356.640 2495.600 358.040 ;
        RECT 4.000 354.640 2498.195 356.640 ;
        RECT 4.400 353.240 2495.600 354.640 ;
        RECT 4.000 351.240 2498.195 353.240 ;
        RECT 4.400 349.840 2495.600 351.240 ;
        RECT 4.000 347.840 2498.195 349.840 ;
        RECT 4.400 346.440 2495.600 347.840 ;
        RECT 4.000 344.440 2498.195 346.440 ;
        RECT 4.400 343.040 2495.600 344.440 ;
        RECT 4.000 341.040 2498.195 343.040 ;
        RECT 4.400 339.640 2495.600 341.040 ;
        RECT 4.000 337.640 2498.195 339.640 ;
        RECT 4.400 336.240 2495.600 337.640 ;
        RECT 4.000 334.240 2498.195 336.240 ;
        RECT 4.400 332.840 2498.195 334.240 ;
        RECT 4.000 330.840 2498.195 332.840 ;
        RECT 4.400 329.440 2495.600 330.840 ;
        RECT 4.000 327.440 2498.195 329.440 ;
        RECT 4.400 326.040 2495.600 327.440 ;
        RECT 4.000 324.040 2498.195 326.040 ;
        RECT 4.000 322.640 2495.600 324.040 ;
        RECT 4.000 320.640 2498.195 322.640 ;
        RECT 4.400 319.240 2495.600 320.640 ;
        RECT 4.000 317.240 2498.195 319.240 ;
        RECT 4.400 315.840 2495.600 317.240 ;
        RECT 4.000 313.840 2498.195 315.840 ;
        RECT 4.400 312.440 2495.600 313.840 ;
        RECT 4.000 310.440 2498.195 312.440 ;
        RECT 4.400 309.040 2495.600 310.440 ;
        RECT 4.000 307.040 2498.195 309.040 ;
        RECT 4.400 305.640 2495.600 307.040 ;
        RECT 4.000 303.640 2498.195 305.640 ;
        RECT 4.400 302.240 2495.600 303.640 ;
        RECT 4.000 300.240 2498.195 302.240 ;
        RECT 4.400 298.840 2495.600 300.240 ;
        RECT 4.000 296.840 2498.195 298.840 ;
        RECT 4.400 295.440 2495.600 296.840 ;
        RECT 4.000 293.440 2498.195 295.440 ;
        RECT 4.400 292.040 2495.600 293.440 ;
        RECT 4.000 290.040 2498.195 292.040 ;
        RECT 4.400 288.640 2495.600 290.040 ;
        RECT 4.000 286.640 2498.195 288.640 ;
        RECT 4.400 285.240 2495.600 286.640 ;
        RECT 4.000 283.240 2498.195 285.240 ;
        RECT 4.400 281.840 2498.195 283.240 ;
        RECT 4.000 279.840 2498.195 281.840 ;
        RECT 4.400 278.440 2495.600 279.840 ;
        RECT 4.000 276.440 2498.195 278.440 ;
        RECT 4.400 275.040 2495.600 276.440 ;
        RECT 4.000 273.040 2498.195 275.040 ;
        RECT 4.400 271.640 2495.600 273.040 ;
        RECT 4.000 269.640 2498.195 271.640 ;
        RECT 4.000 268.240 2495.600 269.640 ;
        RECT 4.000 266.240 2498.195 268.240 ;
        RECT 4.400 264.840 2495.600 266.240 ;
        RECT 4.000 262.840 2498.195 264.840 ;
        RECT 4.400 261.440 2495.600 262.840 ;
        RECT 4.000 259.440 2498.195 261.440 ;
        RECT 4.400 258.040 2495.600 259.440 ;
        RECT 4.000 256.040 2498.195 258.040 ;
        RECT 4.400 254.640 2495.600 256.040 ;
        RECT 4.000 252.640 2498.195 254.640 ;
        RECT 4.400 251.240 2495.600 252.640 ;
        RECT 4.000 249.240 2498.195 251.240 ;
        RECT 4.400 247.840 2495.600 249.240 ;
        RECT 4.000 245.840 2498.195 247.840 ;
        RECT 4.400 244.440 2495.600 245.840 ;
        RECT 4.000 242.440 2498.195 244.440 ;
        RECT 4.400 241.040 2495.600 242.440 ;
        RECT 4.000 239.040 2498.195 241.040 ;
        RECT 4.400 237.640 2495.600 239.040 ;
        RECT 4.000 235.640 2498.195 237.640 ;
        RECT 4.400 234.240 2495.600 235.640 ;
        RECT 4.000 232.240 2498.195 234.240 ;
        RECT 4.400 230.840 2495.600 232.240 ;
        RECT 4.000 228.840 2498.195 230.840 ;
        RECT 4.400 227.440 2498.195 228.840 ;
        RECT 4.000 225.440 2498.195 227.440 ;
        RECT 4.400 224.040 2495.600 225.440 ;
        RECT 4.000 222.040 2498.195 224.040 ;
        RECT 4.400 220.640 2495.600 222.040 ;
        RECT 4.000 218.640 2498.195 220.640 ;
        RECT 4.400 217.240 2495.600 218.640 ;
        RECT 4.000 215.240 2498.195 217.240 ;
        RECT 4.000 213.840 2495.600 215.240 ;
        RECT 4.000 211.840 2498.195 213.840 ;
        RECT 4.400 210.440 2495.600 211.840 ;
        RECT 4.000 208.440 2498.195 210.440 ;
        RECT 4.400 207.040 2495.600 208.440 ;
        RECT 4.000 205.040 2498.195 207.040 ;
        RECT 4.400 203.640 2495.600 205.040 ;
        RECT 4.000 201.640 2498.195 203.640 ;
        RECT 4.400 200.240 2495.600 201.640 ;
        RECT 4.000 198.240 2498.195 200.240 ;
        RECT 4.400 196.840 2495.600 198.240 ;
        RECT 4.000 194.840 2498.195 196.840 ;
        RECT 4.400 193.440 2495.600 194.840 ;
        RECT 4.000 191.440 2498.195 193.440 ;
        RECT 4.400 190.040 2495.600 191.440 ;
        RECT 4.000 188.040 2498.195 190.040 ;
        RECT 4.400 186.640 2495.600 188.040 ;
        RECT 4.000 184.640 2498.195 186.640 ;
        RECT 4.400 183.240 2495.600 184.640 ;
        RECT 4.000 181.240 2498.195 183.240 ;
        RECT 4.400 179.840 2495.600 181.240 ;
        RECT 4.000 177.840 2498.195 179.840 ;
        RECT 4.400 176.440 2495.600 177.840 ;
        RECT 4.000 174.440 2498.195 176.440 ;
        RECT 4.400 173.040 2498.195 174.440 ;
        RECT 4.000 171.040 2498.195 173.040 ;
        RECT 4.400 169.640 2495.600 171.040 ;
        RECT 4.000 167.640 2498.195 169.640 ;
        RECT 4.400 166.240 2495.600 167.640 ;
        RECT 4.000 164.240 2498.195 166.240 ;
        RECT 4.400 162.840 2495.600 164.240 ;
        RECT 4.000 160.840 2498.195 162.840 ;
        RECT 4.000 159.440 2495.600 160.840 ;
        RECT 4.000 157.440 2498.195 159.440 ;
        RECT 4.400 156.040 2495.600 157.440 ;
        RECT 4.000 154.040 2498.195 156.040 ;
        RECT 4.400 152.640 2495.600 154.040 ;
        RECT 4.000 150.640 2498.195 152.640 ;
        RECT 4.400 149.240 2495.600 150.640 ;
        RECT 4.000 147.240 2498.195 149.240 ;
        RECT 4.400 145.840 2495.600 147.240 ;
        RECT 4.000 143.840 2498.195 145.840 ;
        RECT 4.400 142.440 2495.600 143.840 ;
        RECT 4.000 140.440 2498.195 142.440 ;
        RECT 4.400 139.040 2495.600 140.440 ;
        RECT 4.000 137.040 2498.195 139.040 ;
        RECT 4.400 135.640 2495.600 137.040 ;
        RECT 4.000 133.640 2498.195 135.640 ;
        RECT 4.400 132.240 2495.600 133.640 ;
        RECT 4.000 130.240 2498.195 132.240 ;
        RECT 4.400 128.840 2495.600 130.240 ;
        RECT 4.000 126.840 2498.195 128.840 ;
        RECT 4.400 125.440 2495.600 126.840 ;
        RECT 4.000 123.440 2498.195 125.440 ;
        RECT 4.400 122.040 2495.600 123.440 ;
        RECT 4.000 120.040 2498.195 122.040 ;
        RECT 4.400 118.640 2498.195 120.040 ;
        RECT 4.000 116.640 2498.195 118.640 ;
        RECT 4.400 115.240 2495.600 116.640 ;
        RECT 4.000 113.240 2498.195 115.240 ;
        RECT 4.400 111.840 2495.600 113.240 ;
        RECT 4.000 109.840 2498.195 111.840 ;
        RECT 4.400 108.440 2495.600 109.840 ;
        RECT 4.000 106.440 2498.195 108.440 ;
        RECT 4.000 105.040 2495.600 106.440 ;
        RECT 4.000 103.040 2498.195 105.040 ;
        RECT 4.400 101.640 2495.600 103.040 ;
        RECT 4.000 99.640 2498.195 101.640 ;
        RECT 4.400 98.240 2495.600 99.640 ;
        RECT 4.000 96.240 2498.195 98.240 ;
        RECT 4.400 94.840 2495.600 96.240 ;
        RECT 4.000 92.840 2498.195 94.840 ;
        RECT 4.400 91.440 2495.600 92.840 ;
        RECT 4.000 89.440 2498.195 91.440 ;
        RECT 4.400 88.040 2495.600 89.440 ;
        RECT 4.000 86.040 2498.195 88.040 ;
        RECT 4.400 84.640 2495.600 86.040 ;
        RECT 4.000 82.640 2498.195 84.640 ;
        RECT 4.400 81.240 2495.600 82.640 ;
        RECT 4.000 79.240 2498.195 81.240 ;
        RECT 4.400 77.840 2495.600 79.240 ;
        RECT 4.000 75.840 2498.195 77.840 ;
        RECT 4.400 74.440 2495.600 75.840 ;
        RECT 4.000 72.440 2498.195 74.440 ;
        RECT 4.400 71.040 2495.600 72.440 ;
        RECT 4.000 69.040 2498.195 71.040 ;
        RECT 4.400 67.640 2495.600 69.040 ;
        RECT 4.000 65.640 2498.195 67.640 ;
        RECT 4.400 64.240 2498.195 65.640 ;
        RECT 4.000 62.240 2498.195 64.240 ;
        RECT 4.400 60.840 2495.600 62.240 ;
        RECT 4.000 58.840 2498.195 60.840 ;
        RECT 4.400 57.440 2495.600 58.840 ;
        RECT 4.000 55.440 2498.195 57.440 ;
        RECT 4.400 54.040 2495.600 55.440 ;
        RECT 4.000 52.040 2498.195 54.040 ;
        RECT 4.000 50.640 2495.600 52.040 ;
        RECT 4.000 48.640 2498.195 50.640 ;
        RECT 4.400 47.240 2495.600 48.640 ;
        RECT 4.000 45.240 2498.195 47.240 ;
        RECT 4.400 43.840 2495.600 45.240 ;
        RECT 4.000 41.840 2498.195 43.840 ;
        RECT 4.400 40.440 2495.600 41.840 ;
        RECT 4.000 38.440 2498.195 40.440 ;
        RECT 4.400 37.040 2495.600 38.440 ;
        RECT 4.000 35.040 2498.195 37.040 ;
        RECT 4.400 33.640 2495.600 35.040 ;
        RECT 4.000 31.640 2498.195 33.640 ;
        RECT 4.400 30.240 2495.600 31.640 ;
        RECT 4.000 28.240 2498.195 30.240 ;
        RECT 4.400 26.840 2495.600 28.240 ;
        RECT 4.000 24.840 2498.195 26.840 ;
        RECT 4.400 23.440 2495.600 24.840 ;
        RECT 4.000 21.440 2498.195 23.440 ;
        RECT 4.400 20.040 2495.600 21.440 ;
        RECT 4.000 18.040 2498.195 20.040 ;
        RECT 4.400 16.640 2495.600 18.040 ;
        RECT 4.000 14.640 2498.195 16.640 ;
        RECT 4.400 13.240 2495.600 14.640 ;
        RECT 4.000 11.240 2498.195 13.240 ;
        RECT 4.400 9.840 2498.195 11.240 ;
        RECT 4.000 7.840 2498.195 9.840 ;
        RECT 4.400 6.440 2495.600 7.840 ;
        RECT 4.000 4.440 2498.195 6.440 ;
        RECT 4.400 3.040 2495.600 4.440 ;
        RECT 4.000 1.040 2498.195 3.040 ;
        RECT 4.000 0.175 2495.600 1.040 ;
      LAYER met4 ;
        RECT 8.575 2489.440 2492.905 2490.665 ;
        RECT 8.575 10.240 20.640 2489.440 ;
        RECT 23.040 10.240 97.440 2489.440 ;
        RECT 99.840 10.240 174.240 2489.440 ;
        RECT 176.640 10.240 251.040 2489.440 ;
        RECT 253.440 10.240 327.840 2489.440 ;
        RECT 330.240 10.240 404.640 2489.440 ;
        RECT 407.040 10.240 481.440 2489.440 ;
        RECT 483.840 10.240 558.240 2489.440 ;
        RECT 560.640 10.240 635.040 2489.440 ;
        RECT 637.440 10.240 711.840 2489.440 ;
        RECT 714.240 10.240 788.640 2489.440 ;
        RECT 791.040 10.240 865.440 2489.440 ;
        RECT 867.840 10.240 942.240 2489.440 ;
        RECT 944.640 10.240 1019.040 2489.440 ;
        RECT 1021.440 10.240 1095.840 2489.440 ;
        RECT 1098.240 10.240 1172.640 2489.440 ;
        RECT 1175.040 10.240 1249.440 2489.440 ;
        RECT 1251.840 10.240 1326.240 2489.440 ;
        RECT 1328.640 10.240 1403.040 2489.440 ;
        RECT 1405.440 10.240 1479.840 2489.440 ;
        RECT 1482.240 10.240 1556.640 2489.440 ;
        RECT 1559.040 10.240 1633.440 2489.440 ;
        RECT 1635.840 10.240 1710.240 2489.440 ;
        RECT 1712.640 10.240 1787.040 2489.440 ;
        RECT 1789.440 10.240 1863.840 2489.440 ;
        RECT 1866.240 10.240 1940.640 2489.440 ;
        RECT 1943.040 10.240 2017.440 2489.440 ;
        RECT 2019.840 10.240 2094.240 2489.440 ;
        RECT 2096.640 10.240 2171.040 2489.440 ;
        RECT 2173.440 10.240 2247.840 2489.440 ;
        RECT 2250.240 10.240 2324.640 2489.440 ;
        RECT 2327.040 10.240 2401.440 2489.440 ;
        RECT 2403.840 10.240 2478.240 2489.440 ;
        RECT 2480.640 10.240 2492.905 2489.440 ;
        RECT 8.575 6.975 2492.905 10.240 ;
  END
END tile
END LIBRARY


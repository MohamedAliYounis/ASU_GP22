* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for tile abstract view
.subckt tile buffer_processor_data_noc1[0] buffer_processor_data_noc1[10] buffer_processor_data_noc1[11]
+ buffer_processor_data_noc1[12] buffer_processor_data_noc1[13] buffer_processor_data_noc1[14]
+ buffer_processor_data_noc1[15] buffer_processor_data_noc1[16] buffer_processor_data_noc1[17]
+ buffer_processor_data_noc1[18] buffer_processor_data_noc1[19] buffer_processor_data_noc1[1]
+ buffer_processor_data_noc1[20] buffer_processor_data_noc1[21] buffer_processor_data_noc1[22]
+ buffer_processor_data_noc1[23] buffer_processor_data_noc1[24] buffer_processor_data_noc1[25]
+ buffer_processor_data_noc1[26] buffer_processor_data_noc1[27] buffer_processor_data_noc1[28]
+ buffer_processor_data_noc1[29] buffer_processor_data_noc1[2] buffer_processor_data_noc1[30]
+ buffer_processor_data_noc1[31] buffer_processor_data_noc1[32] buffer_processor_data_noc1[33]
+ buffer_processor_data_noc1[34] buffer_processor_data_noc1[35] buffer_processor_data_noc1[36]
+ buffer_processor_data_noc1[37] buffer_processor_data_noc1[38] buffer_processor_data_noc1[39]
+ buffer_processor_data_noc1[3] buffer_processor_data_noc1[40] buffer_processor_data_noc1[41]
+ buffer_processor_data_noc1[42] buffer_processor_data_noc1[43] buffer_processor_data_noc1[44]
+ buffer_processor_data_noc1[45] buffer_processor_data_noc1[46] buffer_processor_data_noc1[47]
+ buffer_processor_data_noc1[48] buffer_processor_data_noc1[49] buffer_processor_data_noc1[4]
+ buffer_processor_data_noc1[50] buffer_processor_data_noc1[51] buffer_processor_data_noc1[52]
+ buffer_processor_data_noc1[53] buffer_processor_data_noc1[54] buffer_processor_data_noc1[55]
+ buffer_processor_data_noc1[56] buffer_processor_data_noc1[57] buffer_processor_data_noc1[58]
+ buffer_processor_data_noc1[59] buffer_processor_data_noc1[5] buffer_processor_data_noc1[60]
+ buffer_processor_data_noc1[61] buffer_processor_data_noc1[62] buffer_processor_data_noc1[63]
+ buffer_processor_data_noc1[6] buffer_processor_data_noc1[7] buffer_processor_data_noc1[8]
+ buffer_processor_data_noc1[9] buffer_processor_data_noc3[0] buffer_processor_data_noc3[10]
+ buffer_processor_data_noc3[11] buffer_processor_data_noc3[12] buffer_processor_data_noc3[13]
+ buffer_processor_data_noc3[14] buffer_processor_data_noc3[15] buffer_processor_data_noc3[16]
+ buffer_processor_data_noc3[17] buffer_processor_data_noc3[18] buffer_processor_data_noc3[19]
+ buffer_processor_data_noc3[1] buffer_processor_data_noc3[20] buffer_processor_data_noc3[21]
+ buffer_processor_data_noc3[22] buffer_processor_data_noc3[23] buffer_processor_data_noc3[24]
+ buffer_processor_data_noc3[25] buffer_processor_data_noc3[26] buffer_processor_data_noc3[27]
+ buffer_processor_data_noc3[28] buffer_processor_data_noc3[29] buffer_processor_data_noc3[2]
+ buffer_processor_data_noc3[30] buffer_processor_data_noc3[31] buffer_processor_data_noc3[32]
+ buffer_processor_data_noc3[33] buffer_processor_data_noc3[34] buffer_processor_data_noc3[35]
+ buffer_processor_data_noc3[36] buffer_processor_data_noc3[37] buffer_processor_data_noc3[38]
+ buffer_processor_data_noc3[39] buffer_processor_data_noc3[3] buffer_processor_data_noc3[40]
+ buffer_processor_data_noc3[41] buffer_processor_data_noc3[42] buffer_processor_data_noc3[43]
+ buffer_processor_data_noc3[44] buffer_processor_data_noc3[45] buffer_processor_data_noc3[46]
+ buffer_processor_data_noc3[47] buffer_processor_data_noc3[48] buffer_processor_data_noc3[49]
+ buffer_processor_data_noc3[4] buffer_processor_data_noc3[50] buffer_processor_data_noc3[51]
+ buffer_processor_data_noc3[52] buffer_processor_data_noc3[53] buffer_processor_data_noc3[54]
+ buffer_processor_data_noc3[55] buffer_processor_data_noc3[56] buffer_processor_data_noc3[57]
+ buffer_processor_data_noc3[58] buffer_processor_data_noc3[59] buffer_processor_data_noc3[5]
+ buffer_processor_data_noc3[60] buffer_processor_data_noc3[61] buffer_processor_data_noc3[62]
+ buffer_processor_data_noc3[63] buffer_processor_data_noc3[6] buffer_processor_data_noc3[7]
+ buffer_processor_data_noc3[8] buffer_processor_data_noc3[9] buffer_processor_valid_noc1
+ buffer_processor_valid_noc3 chipid[0] chipid[10] chipid[11] chipid[12] chipid[13]
+ chipid[1] chipid[2] chipid[3] chipid[4] chipid[5] chipid[6] chipid[7] chipid[8]
+ chipid[9] clk clk_en config_chipid[0] config_chipid[10] config_chipid[11] config_chipid[12]
+ config_chipid[13] config_chipid[1] config_chipid[2] config_chipid[3] config_chipid[4]
+ config_chipid[5] config_chipid[6] config_chipid[7] config_chipid[8] config_chipid[9]
+ config_coreid_x[0] config_coreid_x[1] config_coreid_x[2] config_coreid_x[3] config_coreid_x[4]
+ config_coreid_x[5] config_coreid_x[6] config_coreid_x[7] config_coreid_y[0] config_coreid_y[1]
+ config_coreid_y[2] config_coreid_y[3] config_coreid_y[4] config_coreid_y[5] config_coreid_y[6]
+ config_coreid_y[7] config_csm_en config_hmt_base[0] config_hmt_base[10] config_hmt_base[11]
+ config_hmt_base[12] config_hmt_base[13] config_hmt_base[14] config_hmt_base[15]
+ config_hmt_base[16] config_hmt_base[17] config_hmt_base[18] config_hmt_base[19]
+ config_hmt_base[1] config_hmt_base[20] config_hmt_base[21] config_hmt_base[2] config_hmt_base[3]
+ config_hmt_base[4] config_hmt_base[5] config_hmt_base[6] config_hmt_base[7] config_hmt_base[8]
+ config_hmt_base[9] config_home_alloc_method[0] config_home_alloc_method[1] config_l15_read_res_data_s3[0]
+ config_l15_read_res_data_s3[10] config_l15_read_res_data_s3[11] config_l15_read_res_data_s3[12]
+ config_l15_read_res_data_s3[13] config_l15_read_res_data_s3[14] config_l15_read_res_data_s3[15]
+ config_l15_read_res_data_s3[16] config_l15_read_res_data_s3[17] config_l15_read_res_data_s3[18]
+ config_l15_read_res_data_s3[19] config_l15_read_res_data_s3[1] config_l15_read_res_data_s3[20]
+ config_l15_read_res_data_s3[21] config_l15_read_res_data_s3[22] config_l15_read_res_data_s3[23]
+ config_l15_read_res_data_s3[24] config_l15_read_res_data_s3[25] config_l15_read_res_data_s3[26]
+ config_l15_read_res_data_s3[27] config_l15_read_res_data_s3[28] config_l15_read_res_data_s3[29]
+ config_l15_read_res_data_s3[2] config_l15_read_res_data_s3[30] config_l15_read_res_data_s3[31]
+ config_l15_read_res_data_s3[32] config_l15_read_res_data_s3[33] config_l15_read_res_data_s3[34]
+ config_l15_read_res_data_s3[35] config_l15_read_res_data_s3[36] config_l15_read_res_data_s3[37]
+ config_l15_read_res_data_s3[38] config_l15_read_res_data_s3[39] config_l15_read_res_data_s3[3]
+ config_l15_read_res_data_s3[40] config_l15_read_res_data_s3[41] config_l15_read_res_data_s3[42]
+ config_l15_read_res_data_s3[43] config_l15_read_res_data_s3[44] config_l15_read_res_data_s3[45]
+ config_l15_read_res_data_s3[46] config_l15_read_res_data_s3[47] config_l15_read_res_data_s3[48]
+ config_l15_read_res_data_s3[49] config_l15_read_res_data_s3[4] config_l15_read_res_data_s3[50]
+ config_l15_read_res_data_s3[51] config_l15_read_res_data_s3[52] config_l15_read_res_data_s3[53]
+ config_l15_read_res_data_s3[54] config_l15_read_res_data_s3[55] config_l15_read_res_data_s3[56]
+ config_l15_read_res_data_s3[57] config_l15_read_res_data_s3[58] config_l15_read_res_data_s3[59]
+ config_l15_read_res_data_s3[5] config_l15_read_res_data_s3[60] config_l15_read_res_data_s3[61]
+ config_l15_read_res_data_s3[62] config_l15_read_res_data_s3[63] config_l15_read_res_data_s3[6]
+ config_l15_read_res_data_s3[7] config_l15_read_res_data_s3[8] config_l15_read_res_data_s3[9]
+ config_system_tile_count_5_0[0] config_system_tile_count_5_0[1] config_system_tile_count_5_0[2]
+ config_system_tile_count_5_0[3] config_system_tile_count_5_0[4] config_system_tile_count_5_0[5]
+ coreid_x[0] coreid_x[1] coreid_x[2] coreid_x[3] coreid_x[4] coreid_x[5] coreid_x[6]
+ coreid_x[7] coreid_y[0] coreid_y[1] coreid_y[2] coreid_y[3] coreid_y[4] coreid_y[5]
+ coreid_y[6] coreid_y[7] default_chipid[0] default_chipid[10] default_chipid[11]
+ default_chipid[12] default_chipid[13] default_chipid[1] default_chipid[2] default_chipid[3]
+ default_chipid[4] default_chipid[5] default_chipid[6] default_chipid[7] default_chipid[8]
+ default_chipid[9] default_coreid_x[0] default_coreid_x[1] default_coreid_x[2] default_coreid_x[3]
+ default_coreid_x[4] default_coreid_x[5] default_coreid_x[6] default_coreid_x[7]
+ default_coreid_y[0] default_coreid_y[1] default_coreid_y[2] default_coreid_y[3]
+ default_coreid_y[4] default_coreid_y[5] default_coreid_y[6] default_coreid_y[7]
+ dmbr_l15_stall dummy_core[0] dummy_core[10] dummy_core[11] dummy_core[12] dummy_core[13]
+ dummy_core[14] dummy_core[15] dummy_core[16] dummy_core[17] dummy_core[18] dummy_core[19]
+ dummy_core[1] dummy_core[20] dummy_core[21] dummy_core[22] dummy_core[23] dummy_core[24]
+ dummy_core[25] dummy_core[26] dummy_core[27] dummy_core[28] dummy_core[29] dummy_core[2]
+ dummy_core[30] dummy_core[31] dummy_core[3] dummy_core[4] dummy_core[5] dummy_core[6]
+ dummy_core[7] dummy_core[8] dummy_core[9] dyn0_dEo[0] dyn0_dEo[10] dyn0_dEo[11]
+ dyn0_dEo[12] dyn0_dEo[13] dyn0_dEo[14] dyn0_dEo[15] dyn0_dEo[16] dyn0_dEo[17] dyn0_dEo[18]
+ dyn0_dEo[19] dyn0_dEo[1] dyn0_dEo[20] dyn0_dEo[21] dyn0_dEo[22] dyn0_dEo[23] dyn0_dEo[24]
+ dyn0_dEo[25] dyn0_dEo[26] dyn0_dEo[27] dyn0_dEo[28] dyn0_dEo[29] dyn0_dEo[2] dyn0_dEo[30]
+ dyn0_dEo[31] dyn0_dEo[32] dyn0_dEo[33] dyn0_dEo[34] dyn0_dEo[35] dyn0_dEo[36] dyn0_dEo[37]
+ dyn0_dEo[38] dyn0_dEo[39] dyn0_dEo[3] dyn0_dEo[40] dyn0_dEo[41] dyn0_dEo[42] dyn0_dEo[43]
+ dyn0_dEo[44] dyn0_dEo[45] dyn0_dEo[46] dyn0_dEo[47] dyn0_dEo[48] dyn0_dEo[49] dyn0_dEo[4]
+ dyn0_dEo[50] dyn0_dEo[51] dyn0_dEo[52] dyn0_dEo[53] dyn0_dEo[54] dyn0_dEo[55] dyn0_dEo[56]
+ dyn0_dEo[57] dyn0_dEo[58] dyn0_dEo[59] dyn0_dEo[5] dyn0_dEo[60] dyn0_dEo[61] dyn0_dEo[62]
+ dyn0_dEo[63] dyn0_dEo[6] dyn0_dEo[7] dyn0_dEo[8] dyn0_dEo[9] dyn0_dEo_valid dyn0_dEo_yummy
+ dyn0_dNo[0] dyn0_dNo[10] dyn0_dNo[11] dyn0_dNo[12] dyn0_dNo[13] dyn0_dNo[14] dyn0_dNo[15]
+ dyn0_dNo[16] dyn0_dNo[17] dyn0_dNo[18] dyn0_dNo[19] dyn0_dNo[1] dyn0_dNo[20] dyn0_dNo[21]
+ dyn0_dNo[22] dyn0_dNo[23] dyn0_dNo[24] dyn0_dNo[25] dyn0_dNo[26] dyn0_dNo[27] dyn0_dNo[28]
+ dyn0_dNo[29] dyn0_dNo[2] dyn0_dNo[30] dyn0_dNo[31] dyn0_dNo[32] dyn0_dNo[33] dyn0_dNo[34]
+ dyn0_dNo[35] dyn0_dNo[36] dyn0_dNo[37] dyn0_dNo[38] dyn0_dNo[39] dyn0_dNo[3] dyn0_dNo[40]
+ dyn0_dNo[41] dyn0_dNo[42] dyn0_dNo[43] dyn0_dNo[44] dyn0_dNo[45] dyn0_dNo[46] dyn0_dNo[47]
+ dyn0_dNo[48] dyn0_dNo[49] dyn0_dNo[4] dyn0_dNo[50] dyn0_dNo[51] dyn0_dNo[52] dyn0_dNo[53]
+ dyn0_dNo[54] dyn0_dNo[55] dyn0_dNo[56] dyn0_dNo[57] dyn0_dNo[58] dyn0_dNo[59] dyn0_dNo[5]
+ dyn0_dNo[60] dyn0_dNo[61] dyn0_dNo[62] dyn0_dNo[63] dyn0_dNo[6] dyn0_dNo[7] dyn0_dNo[8]
+ dyn0_dNo[9] dyn0_dNo_valid dyn0_dNo_yummy dyn0_dSo[0] dyn0_dSo[10] dyn0_dSo[11]
+ dyn0_dSo[12] dyn0_dSo[13] dyn0_dSo[14] dyn0_dSo[15] dyn0_dSo[16] dyn0_dSo[17] dyn0_dSo[18]
+ dyn0_dSo[19] dyn0_dSo[1] dyn0_dSo[20] dyn0_dSo[21] dyn0_dSo[22] dyn0_dSo[23] dyn0_dSo[24]
+ dyn0_dSo[25] dyn0_dSo[26] dyn0_dSo[27] dyn0_dSo[28] dyn0_dSo[29] dyn0_dSo[2] dyn0_dSo[30]
+ dyn0_dSo[31] dyn0_dSo[32] dyn0_dSo[33] dyn0_dSo[34] dyn0_dSo[35] dyn0_dSo[36] dyn0_dSo[37]
+ dyn0_dSo[38] dyn0_dSo[39] dyn0_dSo[3] dyn0_dSo[40] dyn0_dSo[41] dyn0_dSo[42] dyn0_dSo[43]
+ dyn0_dSo[44] dyn0_dSo[45] dyn0_dSo[46] dyn0_dSo[47] dyn0_dSo[48] dyn0_dSo[49] dyn0_dSo[4]
+ dyn0_dSo[50] dyn0_dSo[51] dyn0_dSo[52] dyn0_dSo[53] dyn0_dSo[54] dyn0_dSo[55] dyn0_dSo[56]
+ dyn0_dSo[57] dyn0_dSo[58] dyn0_dSo[59] dyn0_dSo[5] dyn0_dSo[60] dyn0_dSo[61] dyn0_dSo[62]
+ dyn0_dSo[63] dyn0_dSo[6] dyn0_dSo[7] dyn0_dSo[8] dyn0_dSo[9] dyn0_dSo_valid dyn0_dSo_yummy
+ dyn0_dWo[0] dyn0_dWo[10] dyn0_dWo[11] dyn0_dWo[12] dyn0_dWo[13] dyn0_dWo[14] dyn0_dWo[15]
+ dyn0_dWo[16] dyn0_dWo[17] dyn0_dWo[18] dyn0_dWo[19] dyn0_dWo[1] dyn0_dWo[20] dyn0_dWo[21]
+ dyn0_dWo[22] dyn0_dWo[23] dyn0_dWo[24] dyn0_dWo[25] dyn0_dWo[26] dyn0_dWo[27] dyn0_dWo[28]
+ dyn0_dWo[29] dyn0_dWo[2] dyn0_dWo[30] dyn0_dWo[31] dyn0_dWo[32] dyn0_dWo[33] dyn0_dWo[34]
+ dyn0_dWo[35] dyn0_dWo[36] dyn0_dWo[37] dyn0_dWo[38] dyn0_dWo[39] dyn0_dWo[3] dyn0_dWo[40]
+ dyn0_dWo[41] dyn0_dWo[42] dyn0_dWo[43] dyn0_dWo[44] dyn0_dWo[45] dyn0_dWo[46] dyn0_dWo[47]
+ dyn0_dWo[48] dyn0_dWo[49] dyn0_dWo[4] dyn0_dWo[50] dyn0_dWo[51] dyn0_dWo[52] dyn0_dWo[53]
+ dyn0_dWo[54] dyn0_dWo[55] dyn0_dWo[56] dyn0_dWo[57] dyn0_dWo[58] dyn0_dWo[59] dyn0_dWo[5]
+ dyn0_dWo[60] dyn0_dWo[61] dyn0_dWo[62] dyn0_dWo[63] dyn0_dWo[6] dyn0_dWo[7] dyn0_dWo[8]
+ dyn0_dWo[9] dyn0_dWo_valid dyn0_dWo_yummy dyn0_dataIn_E[0] dyn0_dataIn_E[10] dyn0_dataIn_E[11]
+ dyn0_dataIn_E[12] dyn0_dataIn_E[13] dyn0_dataIn_E[14] dyn0_dataIn_E[15] dyn0_dataIn_E[16]
+ dyn0_dataIn_E[17] dyn0_dataIn_E[18] dyn0_dataIn_E[19] dyn0_dataIn_E[1] dyn0_dataIn_E[20]
+ dyn0_dataIn_E[21] dyn0_dataIn_E[22] dyn0_dataIn_E[23] dyn0_dataIn_E[24] dyn0_dataIn_E[25]
+ dyn0_dataIn_E[26] dyn0_dataIn_E[27] dyn0_dataIn_E[28] dyn0_dataIn_E[29] dyn0_dataIn_E[2]
+ dyn0_dataIn_E[30] dyn0_dataIn_E[31] dyn0_dataIn_E[32] dyn0_dataIn_E[33] dyn0_dataIn_E[34]
+ dyn0_dataIn_E[35] dyn0_dataIn_E[36] dyn0_dataIn_E[37] dyn0_dataIn_E[38] dyn0_dataIn_E[39]
+ dyn0_dataIn_E[3] dyn0_dataIn_E[40] dyn0_dataIn_E[41] dyn0_dataIn_E[42] dyn0_dataIn_E[43]
+ dyn0_dataIn_E[44] dyn0_dataIn_E[45] dyn0_dataIn_E[46] dyn0_dataIn_E[47] dyn0_dataIn_E[48]
+ dyn0_dataIn_E[49] dyn0_dataIn_E[4] dyn0_dataIn_E[50] dyn0_dataIn_E[51] dyn0_dataIn_E[52]
+ dyn0_dataIn_E[53] dyn0_dataIn_E[54] dyn0_dataIn_E[55] dyn0_dataIn_E[56] dyn0_dataIn_E[57]
+ dyn0_dataIn_E[58] dyn0_dataIn_E[59] dyn0_dataIn_E[5] dyn0_dataIn_E[60] dyn0_dataIn_E[61]
+ dyn0_dataIn_E[62] dyn0_dataIn_E[63] dyn0_dataIn_E[6] dyn0_dataIn_E[7] dyn0_dataIn_E[8]
+ dyn0_dataIn_E[9] dyn0_dataIn_N[0] dyn0_dataIn_N[10] dyn0_dataIn_N[11] dyn0_dataIn_N[12]
+ dyn0_dataIn_N[13] dyn0_dataIn_N[14] dyn0_dataIn_N[15] dyn0_dataIn_N[16] dyn0_dataIn_N[17]
+ dyn0_dataIn_N[18] dyn0_dataIn_N[19] dyn0_dataIn_N[1] dyn0_dataIn_N[20] dyn0_dataIn_N[21]
+ dyn0_dataIn_N[22] dyn0_dataIn_N[23] dyn0_dataIn_N[24] dyn0_dataIn_N[25] dyn0_dataIn_N[26]
+ dyn0_dataIn_N[27] dyn0_dataIn_N[28] dyn0_dataIn_N[29] dyn0_dataIn_N[2] dyn0_dataIn_N[30]
+ dyn0_dataIn_N[31] dyn0_dataIn_N[32] dyn0_dataIn_N[33] dyn0_dataIn_N[34] dyn0_dataIn_N[35]
+ dyn0_dataIn_N[36] dyn0_dataIn_N[37] dyn0_dataIn_N[38] dyn0_dataIn_N[39] dyn0_dataIn_N[3]
+ dyn0_dataIn_N[40] dyn0_dataIn_N[41] dyn0_dataIn_N[42] dyn0_dataIn_N[43] dyn0_dataIn_N[44]
+ dyn0_dataIn_N[45] dyn0_dataIn_N[46] dyn0_dataIn_N[47] dyn0_dataIn_N[48] dyn0_dataIn_N[49]
+ dyn0_dataIn_N[4] dyn0_dataIn_N[50] dyn0_dataIn_N[51] dyn0_dataIn_N[52] dyn0_dataIn_N[53]
+ dyn0_dataIn_N[54] dyn0_dataIn_N[55] dyn0_dataIn_N[56] dyn0_dataIn_N[57] dyn0_dataIn_N[58]
+ dyn0_dataIn_N[59] dyn0_dataIn_N[5] dyn0_dataIn_N[60] dyn0_dataIn_N[61] dyn0_dataIn_N[62]
+ dyn0_dataIn_N[63] dyn0_dataIn_N[6] dyn0_dataIn_N[7] dyn0_dataIn_N[8] dyn0_dataIn_N[9]
+ dyn0_dataIn_S[0] dyn0_dataIn_S[10] dyn0_dataIn_S[11] dyn0_dataIn_S[12] dyn0_dataIn_S[13]
+ dyn0_dataIn_S[14] dyn0_dataIn_S[15] dyn0_dataIn_S[16] dyn0_dataIn_S[17] dyn0_dataIn_S[18]
+ dyn0_dataIn_S[19] dyn0_dataIn_S[1] dyn0_dataIn_S[20] dyn0_dataIn_S[21] dyn0_dataIn_S[22]
+ dyn0_dataIn_S[23] dyn0_dataIn_S[24] dyn0_dataIn_S[25] dyn0_dataIn_S[26] dyn0_dataIn_S[27]
+ dyn0_dataIn_S[28] dyn0_dataIn_S[29] dyn0_dataIn_S[2] dyn0_dataIn_S[30] dyn0_dataIn_S[31]
+ dyn0_dataIn_S[32] dyn0_dataIn_S[33] dyn0_dataIn_S[34] dyn0_dataIn_S[35] dyn0_dataIn_S[36]
+ dyn0_dataIn_S[37] dyn0_dataIn_S[38] dyn0_dataIn_S[39] dyn0_dataIn_S[3] dyn0_dataIn_S[40]
+ dyn0_dataIn_S[41] dyn0_dataIn_S[42] dyn0_dataIn_S[43] dyn0_dataIn_S[44] dyn0_dataIn_S[45]
+ dyn0_dataIn_S[46] dyn0_dataIn_S[47] dyn0_dataIn_S[48] dyn0_dataIn_S[49] dyn0_dataIn_S[4]
+ dyn0_dataIn_S[50] dyn0_dataIn_S[51] dyn0_dataIn_S[52] dyn0_dataIn_S[53] dyn0_dataIn_S[54]
+ dyn0_dataIn_S[55] dyn0_dataIn_S[56] dyn0_dataIn_S[57] dyn0_dataIn_S[58] dyn0_dataIn_S[59]
+ dyn0_dataIn_S[5] dyn0_dataIn_S[60] dyn0_dataIn_S[61] dyn0_dataIn_S[62] dyn0_dataIn_S[63]
+ dyn0_dataIn_S[6] dyn0_dataIn_S[7] dyn0_dataIn_S[8] dyn0_dataIn_S[9] dyn0_dataIn_W[0]
+ dyn0_dataIn_W[10] dyn0_dataIn_W[11] dyn0_dataIn_W[12] dyn0_dataIn_W[13] dyn0_dataIn_W[14]
+ dyn0_dataIn_W[15] dyn0_dataIn_W[16] dyn0_dataIn_W[17] dyn0_dataIn_W[18] dyn0_dataIn_W[19]
+ dyn0_dataIn_W[1] dyn0_dataIn_W[20] dyn0_dataIn_W[21] dyn0_dataIn_W[22] dyn0_dataIn_W[23]
+ dyn0_dataIn_W[24] dyn0_dataIn_W[25] dyn0_dataIn_W[26] dyn0_dataIn_W[27] dyn0_dataIn_W[28]
+ dyn0_dataIn_W[29] dyn0_dataIn_W[2] dyn0_dataIn_W[30] dyn0_dataIn_W[31] dyn0_dataIn_W[32]
+ dyn0_dataIn_W[33] dyn0_dataIn_W[34] dyn0_dataIn_W[35] dyn0_dataIn_W[36] dyn0_dataIn_W[37]
+ dyn0_dataIn_W[38] dyn0_dataIn_W[39] dyn0_dataIn_W[3] dyn0_dataIn_W[40] dyn0_dataIn_W[41]
+ dyn0_dataIn_W[42] dyn0_dataIn_W[43] dyn0_dataIn_W[44] dyn0_dataIn_W[45] dyn0_dataIn_W[46]
+ dyn0_dataIn_W[47] dyn0_dataIn_W[48] dyn0_dataIn_W[49] dyn0_dataIn_W[4] dyn0_dataIn_W[50]
+ dyn0_dataIn_W[51] dyn0_dataIn_W[52] dyn0_dataIn_W[53] dyn0_dataIn_W[54] dyn0_dataIn_W[55]
+ dyn0_dataIn_W[56] dyn0_dataIn_W[57] dyn0_dataIn_W[58] dyn0_dataIn_W[59] dyn0_dataIn_W[5]
+ dyn0_dataIn_W[60] dyn0_dataIn_W[61] dyn0_dataIn_W[62] dyn0_dataIn_W[63] dyn0_dataIn_W[6]
+ dyn0_dataIn_W[7] dyn0_dataIn_W[8] dyn0_dataIn_W[9] dyn0_validIn_E dyn0_validIn_N
+ dyn0_validIn_S dyn0_validIn_W dyn0_yummyOut_E dyn0_yummyOut_N dyn0_yummyOut_S dyn0_yummyOut_W
+ dyn1_dEo[0] dyn1_dEo[10] dyn1_dEo[11] dyn1_dEo[12] dyn1_dEo[13] dyn1_dEo[14] dyn1_dEo[15]
+ dyn1_dEo[16] dyn1_dEo[17] dyn1_dEo[18] dyn1_dEo[19] dyn1_dEo[1] dyn1_dEo[20] dyn1_dEo[21]
+ dyn1_dEo[22] dyn1_dEo[23] dyn1_dEo[24] dyn1_dEo[25] dyn1_dEo[26] dyn1_dEo[27] dyn1_dEo[28]
+ dyn1_dEo[29] dyn1_dEo[2] dyn1_dEo[30] dyn1_dEo[31] dyn1_dEo[32] dyn1_dEo[33] dyn1_dEo[34]
+ dyn1_dEo[35] dyn1_dEo[36] dyn1_dEo[37] dyn1_dEo[38] dyn1_dEo[39] dyn1_dEo[3] dyn1_dEo[40]
+ dyn1_dEo[41] dyn1_dEo[42] dyn1_dEo[43] dyn1_dEo[44] dyn1_dEo[45] dyn1_dEo[46] dyn1_dEo[47]
+ dyn1_dEo[48] dyn1_dEo[49] dyn1_dEo[4] dyn1_dEo[50] dyn1_dEo[51] dyn1_dEo[52] dyn1_dEo[53]
+ dyn1_dEo[54] dyn1_dEo[55] dyn1_dEo[56] dyn1_dEo[57] dyn1_dEo[58] dyn1_dEo[59] dyn1_dEo[5]
+ dyn1_dEo[60] dyn1_dEo[61] dyn1_dEo[62] dyn1_dEo[63] dyn1_dEo[6] dyn1_dEo[7] dyn1_dEo[8]
+ dyn1_dEo[9] dyn1_dEo_valid dyn1_dEo_yummy dyn1_dNo[0] dyn1_dNo[10] dyn1_dNo[11]
+ dyn1_dNo[12] dyn1_dNo[13] dyn1_dNo[14] dyn1_dNo[15] dyn1_dNo[16] dyn1_dNo[17] dyn1_dNo[18]
+ dyn1_dNo[19] dyn1_dNo[1] dyn1_dNo[20] dyn1_dNo[21] dyn1_dNo[22] dyn1_dNo[23] dyn1_dNo[24]
+ dyn1_dNo[25] dyn1_dNo[26] dyn1_dNo[27] dyn1_dNo[28] dyn1_dNo[29] dyn1_dNo[2] dyn1_dNo[30]
+ dyn1_dNo[31] dyn1_dNo[32] dyn1_dNo[33] dyn1_dNo[34] dyn1_dNo[35] dyn1_dNo[36] dyn1_dNo[37]
+ dyn1_dNo[38] dyn1_dNo[39] dyn1_dNo[3] dyn1_dNo[40] dyn1_dNo[41] dyn1_dNo[42] dyn1_dNo[43]
+ dyn1_dNo[44] dyn1_dNo[45] dyn1_dNo[46] dyn1_dNo[47] dyn1_dNo[48] dyn1_dNo[49] dyn1_dNo[4]
+ dyn1_dNo[50] dyn1_dNo[51] dyn1_dNo[52] dyn1_dNo[53] dyn1_dNo[54] dyn1_dNo[55] dyn1_dNo[56]
+ dyn1_dNo[57] dyn1_dNo[58] dyn1_dNo[59] dyn1_dNo[5] dyn1_dNo[60] dyn1_dNo[61] dyn1_dNo[62]
+ dyn1_dNo[63] dyn1_dNo[6] dyn1_dNo[7] dyn1_dNo[8] dyn1_dNo[9] dyn1_dNo_valid dyn1_dNo_yummy
+ dyn1_dSo[0] dyn1_dSo[10] dyn1_dSo[11] dyn1_dSo[12] dyn1_dSo[13] dyn1_dSo[14] dyn1_dSo[15]
+ dyn1_dSo[16] dyn1_dSo[17] dyn1_dSo[18] dyn1_dSo[19] dyn1_dSo[1] dyn1_dSo[20] dyn1_dSo[21]
+ dyn1_dSo[22] dyn1_dSo[23] dyn1_dSo[24] dyn1_dSo[25] dyn1_dSo[26] dyn1_dSo[27] dyn1_dSo[28]
+ dyn1_dSo[29] dyn1_dSo[2] dyn1_dSo[30] dyn1_dSo[31] dyn1_dSo[32] dyn1_dSo[33] dyn1_dSo[34]
+ dyn1_dSo[35] dyn1_dSo[36] dyn1_dSo[37] dyn1_dSo[38] dyn1_dSo[39] dyn1_dSo[3] dyn1_dSo[40]
+ dyn1_dSo[41] dyn1_dSo[42] dyn1_dSo[43] dyn1_dSo[44] dyn1_dSo[45] dyn1_dSo[46] dyn1_dSo[47]
+ dyn1_dSo[48] dyn1_dSo[49] dyn1_dSo[4] dyn1_dSo[50] dyn1_dSo[51] dyn1_dSo[52] dyn1_dSo[53]
+ dyn1_dSo[54] dyn1_dSo[55] dyn1_dSo[56] dyn1_dSo[57] dyn1_dSo[58] dyn1_dSo[59] dyn1_dSo[5]
+ dyn1_dSo[60] dyn1_dSo[61] dyn1_dSo[62] dyn1_dSo[63] dyn1_dSo[6] dyn1_dSo[7] dyn1_dSo[8]
+ dyn1_dSo[9] dyn1_dSo_valid dyn1_dSo_yummy dyn1_dWo[0] dyn1_dWo[10] dyn1_dWo[11]
+ dyn1_dWo[12] dyn1_dWo[13] dyn1_dWo[14] dyn1_dWo[15] dyn1_dWo[16] dyn1_dWo[17] dyn1_dWo[18]
+ dyn1_dWo[19] dyn1_dWo[1] dyn1_dWo[20] dyn1_dWo[21] dyn1_dWo[22] dyn1_dWo[23] dyn1_dWo[24]
+ dyn1_dWo[25] dyn1_dWo[26] dyn1_dWo[27] dyn1_dWo[28] dyn1_dWo[29] dyn1_dWo[2] dyn1_dWo[30]
+ dyn1_dWo[31] dyn1_dWo[32] dyn1_dWo[33] dyn1_dWo[34] dyn1_dWo[35] dyn1_dWo[36] dyn1_dWo[37]
+ dyn1_dWo[38] dyn1_dWo[39] dyn1_dWo[3] dyn1_dWo[40] dyn1_dWo[41] dyn1_dWo[42] dyn1_dWo[43]
+ dyn1_dWo[44] dyn1_dWo[45] dyn1_dWo[46] dyn1_dWo[47] dyn1_dWo[48] dyn1_dWo[49] dyn1_dWo[4]
+ dyn1_dWo[50] dyn1_dWo[51] dyn1_dWo[52] dyn1_dWo[53] dyn1_dWo[54] dyn1_dWo[55] dyn1_dWo[56]
+ dyn1_dWo[57] dyn1_dWo[58] dyn1_dWo[59] dyn1_dWo[5] dyn1_dWo[60] dyn1_dWo[61] dyn1_dWo[62]
+ dyn1_dWo[63] dyn1_dWo[6] dyn1_dWo[7] dyn1_dWo[8] dyn1_dWo[9] dyn1_dWo_valid dyn1_dWo_yummy
+ dyn1_dataIn_E[0] dyn1_dataIn_E[10] dyn1_dataIn_E[11] dyn1_dataIn_E[12] dyn1_dataIn_E[13]
+ dyn1_dataIn_E[14] dyn1_dataIn_E[15] dyn1_dataIn_E[16] dyn1_dataIn_E[17] dyn1_dataIn_E[18]
+ dyn1_dataIn_E[19] dyn1_dataIn_E[1] dyn1_dataIn_E[20] dyn1_dataIn_E[21] dyn1_dataIn_E[22]
+ dyn1_dataIn_E[23] dyn1_dataIn_E[24] dyn1_dataIn_E[25] dyn1_dataIn_E[26] dyn1_dataIn_E[27]
+ dyn1_dataIn_E[28] dyn1_dataIn_E[29] dyn1_dataIn_E[2] dyn1_dataIn_E[30] dyn1_dataIn_E[31]
+ dyn1_dataIn_E[32] dyn1_dataIn_E[33] dyn1_dataIn_E[34] dyn1_dataIn_E[35] dyn1_dataIn_E[36]
+ dyn1_dataIn_E[37] dyn1_dataIn_E[38] dyn1_dataIn_E[39] dyn1_dataIn_E[3] dyn1_dataIn_E[40]
+ dyn1_dataIn_E[41] dyn1_dataIn_E[42] dyn1_dataIn_E[43] dyn1_dataIn_E[44] dyn1_dataIn_E[45]
+ dyn1_dataIn_E[46] dyn1_dataIn_E[47] dyn1_dataIn_E[48] dyn1_dataIn_E[49] dyn1_dataIn_E[4]
+ dyn1_dataIn_E[50] dyn1_dataIn_E[51] dyn1_dataIn_E[52] dyn1_dataIn_E[53] dyn1_dataIn_E[54]
+ dyn1_dataIn_E[55] dyn1_dataIn_E[56] dyn1_dataIn_E[57] dyn1_dataIn_E[58] dyn1_dataIn_E[59]
+ dyn1_dataIn_E[5] dyn1_dataIn_E[60] dyn1_dataIn_E[61] dyn1_dataIn_E[62] dyn1_dataIn_E[63]
+ dyn1_dataIn_E[6] dyn1_dataIn_E[7] dyn1_dataIn_E[8] dyn1_dataIn_E[9] dyn1_dataIn_N[0]
+ dyn1_dataIn_N[10] dyn1_dataIn_N[11] dyn1_dataIn_N[12] dyn1_dataIn_N[13] dyn1_dataIn_N[14]
+ dyn1_dataIn_N[15] dyn1_dataIn_N[16] dyn1_dataIn_N[17] dyn1_dataIn_N[18] dyn1_dataIn_N[19]
+ dyn1_dataIn_N[1] dyn1_dataIn_N[20] dyn1_dataIn_N[21] dyn1_dataIn_N[22] dyn1_dataIn_N[23]
+ dyn1_dataIn_N[24] dyn1_dataIn_N[25] dyn1_dataIn_N[26] dyn1_dataIn_N[27] dyn1_dataIn_N[28]
+ dyn1_dataIn_N[29] dyn1_dataIn_N[2] dyn1_dataIn_N[30] dyn1_dataIn_N[31] dyn1_dataIn_N[32]
+ dyn1_dataIn_N[33] dyn1_dataIn_N[34] dyn1_dataIn_N[35] dyn1_dataIn_N[36] dyn1_dataIn_N[37]
+ dyn1_dataIn_N[38] dyn1_dataIn_N[39] dyn1_dataIn_N[3] dyn1_dataIn_N[40] dyn1_dataIn_N[41]
+ dyn1_dataIn_N[42] dyn1_dataIn_N[43] dyn1_dataIn_N[44] dyn1_dataIn_N[45] dyn1_dataIn_N[46]
+ dyn1_dataIn_N[47] dyn1_dataIn_N[48] dyn1_dataIn_N[49] dyn1_dataIn_N[4] dyn1_dataIn_N[50]
+ dyn1_dataIn_N[51] dyn1_dataIn_N[52] dyn1_dataIn_N[53] dyn1_dataIn_N[54] dyn1_dataIn_N[55]
+ dyn1_dataIn_N[56] dyn1_dataIn_N[57] dyn1_dataIn_N[58] dyn1_dataIn_N[59] dyn1_dataIn_N[5]
+ dyn1_dataIn_N[60] dyn1_dataIn_N[61] dyn1_dataIn_N[62] dyn1_dataIn_N[63] dyn1_dataIn_N[6]
+ dyn1_dataIn_N[7] dyn1_dataIn_N[8] dyn1_dataIn_N[9] dyn1_dataIn_S[0] dyn1_dataIn_S[10]
+ dyn1_dataIn_S[11] dyn1_dataIn_S[12] dyn1_dataIn_S[13] dyn1_dataIn_S[14] dyn1_dataIn_S[15]
+ dyn1_dataIn_S[16] dyn1_dataIn_S[17] dyn1_dataIn_S[18] dyn1_dataIn_S[19] dyn1_dataIn_S[1]
+ dyn1_dataIn_S[20] dyn1_dataIn_S[21] dyn1_dataIn_S[22] dyn1_dataIn_S[23] dyn1_dataIn_S[24]
+ dyn1_dataIn_S[25] dyn1_dataIn_S[26] dyn1_dataIn_S[27] dyn1_dataIn_S[28] dyn1_dataIn_S[29]
+ dyn1_dataIn_S[2] dyn1_dataIn_S[30] dyn1_dataIn_S[31] dyn1_dataIn_S[32] dyn1_dataIn_S[33]
+ dyn1_dataIn_S[34] dyn1_dataIn_S[35] dyn1_dataIn_S[36] dyn1_dataIn_S[37] dyn1_dataIn_S[38]
+ dyn1_dataIn_S[39] dyn1_dataIn_S[3] dyn1_dataIn_S[40] dyn1_dataIn_S[41] dyn1_dataIn_S[42]
+ dyn1_dataIn_S[43] dyn1_dataIn_S[44] dyn1_dataIn_S[45] dyn1_dataIn_S[46] dyn1_dataIn_S[47]
+ dyn1_dataIn_S[48] dyn1_dataIn_S[49] dyn1_dataIn_S[4] dyn1_dataIn_S[50] dyn1_dataIn_S[51]
+ dyn1_dataIn_S[52] dyn1_dataIn_S[53] dyn1_dataIn_S[54] dyn1_dataIn_S[55] dyn1_dataIn_S[56]
+ dyn1_dataIn_S[57] dyn1_dataIn_S[58] dyn1_dataIn_S[59] dyn1_dataIn_S[5] dyn1_dataIn_S[60]
+ dyn1_dataIn_S[61] dyn1_dataIn_S[62] dyn1_dataIn_S[63] dyn1_dataIn_S[6] dyn1_dataIn_S[7]
+ dyn1_dataIn_S[8] dyn1_dataIn_S[9] dyn1_dataIn_W[0] dyn1_dataIn_W[10] dyn1_dataIn_W[11]
+ dyn1_dataIn_W[12] dyn1_dataIn_W[13] dyn1_dataIn_W[14] dyn1_dataIn_W[15] dyn1_dataIn_W[16]
+ dyn1_dataIn_W[17] dyn1_dataIn_W[18] dyn1_dataIn_W[19] dyn1_dataIn_W[1] dyn1_dataIn_W[20]
+ dyn1_dataIn_W[21] dyn1_dataIn_W[22] dyn1_dataIn_W[23] dyn1_dataIn_W[24] dyn1_dataIn_W[25]
+ dyn1_dataIn_W[26] dyn1_dataIn_W[27] dyn1_dataIn_W[28] dyn1_dataIn_W[29] dyn1_dataIn_W[2]
+ dyn1_dataIn_W[30] dyn1_dataIn_W[31] dyn1_dataIn_W[32] dyn1_dataIn_W[33] dyn1_dataIn_W[34]
+ dyn1_dataIn_W[35] dyn1_dataIn_W[36] dyn1_dataIn_W[37] dyn1_dataIn_W[38] dyn1_dataIn_W[39]
+ dyn1_dataIn_W[3] dyn1_dataIn_W[40] dyn1_dataIn_W[41] dyn1_dataIn_W[42] dyn1_dataIn_W[43]
+ dyn1_dataIn_W[44] dyn1_dataIn_W[45] dyn1_dataIn_W[46] dyn1_dataIn_W[47] dyn1_dataIn_W[48]
+ dyn1_dataIn_W[49] dyn1_dataIn_W[4] dyn1_dataIn_W[50] dyn1_dataIn_W[51] dyn1_dataIn_W[52]
+ dyn1_dataIn_W[53] dyn1_dataIn_W[54] dyn1_dataIn_W[55] dyn1_dataIn_W[56] dyn1_dataIn_W[57]
+ dyn1_dataIn_W[58] dyn1_dataIn_W[59] dyn1_dataIn_W[5] dyn1_dataIn_W[60] dyn1_dataIn_W[61]
+ dyn1_dataIn_W[62] dyn1_dataIn_W[63] dyn1_dataIn_W[6] dyn1_dataIn_W[7] dyn1_dataIn_W[8]
+ dyn1_dataIn_W[9] dyn1_validIn_E dyn1_validIn_N dyn1_validIn_S dyn1_validIn_W dyn1_yummyOut_E
+ dyn1_yummyOut_N dyn1_yummyOut_S dyn1_yummyOut_W dyn2_dEo[0] dyn2_dEo[10] dyn2_dEo[11]
+ dyn2_dEo[12] dyn2_dEo[13] dyn2_dEo[14] dyn2_dEo[15] dyn2_dEo[16] dyn2_dEo[17] dyn2_dEo[18]
+ dyn2_dEo[19] dyn2_dEo[1] dyn2_dEo[20] dyn2_dEo[21] dyn2_dEo[22] dyn2_dEo[23] dyn2_dEo[24]
+ dyn2_dEo[25] dyn2_dEo[26] dyn2_dEo[27] dyn2_dEo[28] dyn2_dEo[29] dyn2_dEo[2] dyn2_dEo[30]
+ dyn2_dEo[31] dyn2_dEo[32] dyn2_dEo[33] dyn2_dEo[34] dyn2_dEo[35] dyn2_dEo[36] dyn2_dEo[37]
+ dyn2_dEo[38] dyn2_dEo[39] dyn2_dEo[3] dyn2_dEo[40] dyn2_dEo[41] dyn2_dEo[42] dyn2_dEo[43]
+ dyn2_dEo[44] dyn2_dEo[45] dyn2_dEo[46] dyn2_dEo[47] dyn2_dEo[48] dyn2_dEo[49] dyn2_dEo[4]
+ dyn2_dEo[50] dyn2_dEo[51] dyn2_dEo[52] dyn2_dEo[53] dyn2_dEo[54] dyn2_dEo[55] dyn2_dEo[56]
+ dyn2_dEo[57] dyn2_dEo[58] dyn2_dEo[59] dyn2_dEo[5] dyn2_dEo[60] dyn2_dEo[61] dyn2_dEo[62]
+ dyn2_dEo[63] dyn2_dEo[6] dyn2_dEo[7] dyn2_dEo[8] dyn2_dEo[9] dyn2_dEo_valid dyn2_dEo_yummy
+ dyn2_dNo[0] dyn2_dNo[10] dyn2_dNo[11] dyn2_dNo[12] dyn2_dNo[13] dyn2_dNo[14] dyn2_dNo[15]
+ dyn2_dNo[16] dyn2_dNo[17] dyn2_dNo[18] dyn2_dNo[19] dyn2_dNo[1] dyn2_dNo[20] dyn2_dNo[21]
+ dyn2_dNo[22] dyn2_dNo[23] dyn2_dNo[24] dyn2_dNo[25] dyn2_dNo[26] dyn2_dNo[27] dyn2_dNo[28]
+ dyn2_dNo[29] dyn2_dNo[2] dyn2_dNo[30] dyn2_dNo[31] dyn2_dNo[32] dyn2_dNo[33] dyn2_dNo[34]
+ dyn2_dNo[35] dyn2_dNo[36] dyn2_dNo[37] dyn2_dNo[38] dyn2_dNo[39] dyn2_dNo[3] dyn2_dNo[40]
+ dyn2_dNo[41] dyn2_dNo[42] dyn2_dNo[43] dyn2_dNo[44] dyn2_dNo[45] dyn2_dNo[46] dyn2_dNo[47]
+ dyn2_dNo[48] dyn2_dNo[49] dyn2_dNo[4] dyn2_dNo[50] dyn2_dNo[51] dyn2_dNo[52] dyn2_dNo[53]
+ dyn2_dNo[54] dyn2_dNo[55] dyn2_dNo[56] dyn2_dNo[57] dyn2_dNo[58] dyn2_dNo[59] dyn2_dNo[5]
+ dyn2_dNo[60] dyn2_dNo[61] dyn2_dNo[62] dyn2_dNo[63] dyn2_dNo[6] dyn2_dNo[7] dyn2_dNo[8]
+ dyn2_dNo[9] dyn2_dNo_valid dyn2_dNo_yummy dyn2_dSo[0] dyn2_dSo[10] dyn2_dSo[11]
+ dyn2_dSo[12] dyn2_dSo[13] dyn2_dSo[14] dyn2_dSo[15] dyn2_dSo[16] dyn2_dSo[17] dyn2_dSo[18]
+ dyn2_dSo[19] dyn2_dSo[1] dyn2_dSo[20] dyn2_dSo[21] dyn2_dSo[22] dyn2_dSo[23] dyn2_dSo[24]
+ dyn2_dSo[25] dyn2_dSo[26] dyn2_dSo[27] dyn2_dSo[28] dyn2_dSo[29] dyn2_dSo[2] dyn2_dSo[30]
+ dyn2_dSo[31] dyn2_dSo[32] dyn2_dSo[33] dyn2_dSo[34] dyn2_dSo[35] dyn2_dSo[36] dyn2_dSo[37]
+ dyn2_dSo[38] dyn2_dSo[39] dyn2_dSo[3] dyn2_dSo[40] dyn2_dSo[41] dyn2_dSo[42] dyn2_dSo[43]
+ dyn2_dSo[44] dyn2_dSo[45] dyn2_dSo[46] dyn2_dSo[47] dyn2_dSo[48] dyn2_dSo[49] dyn2_dSo[4]
+ dyn2_dSo[50] dyn2_dSo[51] dyn2_dSo[52] dyn2_dSo[53] dyn2_dSo[54] dyn2_dSo[55] dyn2_dSo[56]
+ dyn2_dSo[57] dyn2_dSo[58] dyn2_dSo[59] dyn2_dSo[5] dyn2_dSo[60] dyn2_dSo[61] dyn2_dSo[62]
+ dyn2_dSo[63] dyn2_dSo[6] dyn2_dSo[7] dyn2_dSo[8] dyn2_dSo[9] dyn2_dSo_valid dyn2_dSo_yummy
+ dyn2_dWo[0] dyn2_dWo[10] dyn2_dWo[11] dyn2_dWo[12] dyn2_dWo[13] dyn2_dWo[14] dyn2_dWo[15]
+ dyn2_dWo[16] dyn2_dWo[17] dyn2_dWo[18] dyn2_dWo[19] dyn2_dWo[1] dyn2_dWo[20] dyn2_dWo[21]
+ dyn2_dWo[22] dyn2_dWo[23] dyn2_dWo[24] dyn2_dWo[25] dyn2_dWo[26] dyn2_dWo[27] dyn2_dWo[28]
+ dyn2_dWo[29] dyn2_dWo[2] dyn2_dWo[30] dyn2_dWo[31] dyn2_dWo[32] dyn2_dWo[33] dyn2_dWo[34]
+ dyn2_dWo[35] dyn2_dWo[36] dyn2_dWo[37] dyn2_dWo[38] dyn2_dWo[39] dyn2_dWo[3] dyn2_dWo[40]
+ dyn2_dWo[41] dyn2_dWo[42] dyn2_dWo[43] dyn2_dWo[44] dyn2_dWo[45] dyn2_dWo[46] dyn2_dWo[47]
+ dyn2_dWo[48] dyn2_dWo[49] dyn2_dWo[4] dyn2_dWo[50] dyn2_dWo[51] dyn2_dWo[52] dyn2_dWo[53]
+ dyn2_dWo[54] dyn2_dWo[55] dyn2_dWo[56] dyn2_dWo[57] dyn2_dWo[58] dyn2_dWo[59] dyn2_dWo[5]
+ dyn2_dWo[60] dyn2_dWo[61] dyn2_dWo[62] dyn2_dWo[63] dyn2_dWo[6] dyn2_dWo[7] dyn2_dWo[8]
+ dyn2_dWo[9] dyn2_dWo_valid dyn2_dWo_yummy dyn2_dataIn_E[0] dyn2_dataIn_E[10] dyn2_dataIn_E[11]
+ dyn2_dataIn_E[12] dyn2_dataIn_E[13] dyn2_dataIn_E[14] dyn2_dataIn_E[15] dyn2_dataIn_E[16]
+ dyn2_dataIn_E[17] dyn2_dataIn_E[18] dyn2_dataIn_E[19] dyn2_dataIn_E[1] dyn2_dataIn_E[20]
+ dyn2_dataIn_E[21] dyn2_dataIn_E[22] dyn2_dataIn_E[23] dyn2_dataIn_E[24] dyn2_dataIn_E[25]
+ dyn2_dataIn_E[26] dyn2_dataIn_E[27] dyn2_dataIn_E[28] dyn2_dataIn_E[29] dyn2_dataIn_E[2]
+ dyn2_dataIn_E[30] dyn2_dataIn_E[31] dyn2_dataIn_E[32] dyn2_dataIn_E[33] dyn2_dataIn_E[34]
+ dyn2_dataIn_E[35] dyn2_dataIn_E[36] dyn2_dataIn_E[37] dyn2_dataIn_E[38] dyn2_dataIn_E[39]
+ dyn2_dataIn_E[3] dyn2_dataIn_E[40] dyn2_dataIn_E[41] dyn2_dataIn_E[42] dyn2_dataIn_E[43]
+ dyn2_dataIn_E[44] dyn2_dataIn_E[45] dyn2_dataIn_E[46] dyn2_dataIn_E[47] dyn2_dataIn_E[48]
+ dyn2_dataIn_E[49] dyn2_dataIn_E[4] dyn2_dataIn_E[50] dyn2_dataIn_E[51] dyn2_dataIn_E[52]
+ dyn2_dataIn_E[53] dyn2_dataIn_E[54] dyn2_dataIn_E[55] dyn2_dataIn_E[56] dyn2_dataIn_E[57]
+ dyn2_dataIn_E[58] dyn2_dataIn_E[59] dyn2_dataIn_E[5] dyn2_dataIn_E[60] dyn2_dataIn_E[61]
+ dyn2_dataIn_E[62] dyn2_dataIn_E[63] dyn2_dataIn_E[6] dyn2_dataIn_E[7] dyn2_dataIn_E[8]
+ dyn2_dataIn_E[9] dyn2_dataIn_N[0] dyn2_dataIn_N[10] dyn2_dataIn_N[11] dyn2_dataIn_N[12]
+ dyn2_dataIn_N[13] dyn2_dataIn_N[14] dyn2_dataIn_N[15] dyn2_dataIn_N[16] dyn2_dataIn_N[17]
+ dyn2_dataIn_N[18] dyn2_dataIn_N[19] dyn2_dataIn_N[1] dyn2_dataIn_N[20] dyn2_dataIn_N[21]
+ dyn2_dataIn_N[22] dyn2_dataIn_N[23] dyn2_dataIn_N[24] dyn2_dataIn_N[25] dyn2_dataIn_N[26]
+ dyn2_dataIn_N[27] dyn2_dataIn_N[28] dyn2_dataIn_N[29] dyn2_dataIn_N[2] dyn2_dataIn_N[30]
+ dyn2_dataIn_N[31] dyn2_dataIn_N[32] dyn2_dataIn_N[33] dyn2_dataIn_N[34] dyn2_dataIn_N[35]
+ dyn2_dataIn_N[36] dyn2_dataIn_N[37] dyn2_dataIn_N[38] dyn2_dataIn_N[39] dyn2_dataIn_N[3]
+ dyn2_dataIn_N[40] dyn2_dataIn_N[41] dyn2_dataIn_N[42] dyn2_dataIn_N[43] dyn2_dataIn_N[44]
+ dyn2_dataIn_N[45] dyn2_dataIn_N[46] dyn2_dataIn_N[47] dyn2_dataIn_N[48] dyn2_dataIn_N[49]
+ dyn2_dataIn_N[4] dyn2_dataIn_N[50] dyn2_dataIn_N[51] dyn2_dataIn_N[52] dyn2_dataIn_N[53]
+ dyn2_dataIn_N[54] dyn2_dataIn_N[55] dyn2_dataIn_N[56] dyn2_dataIn_N[57] dyn2_dataIn_N[58]
+ dyn2_dataIn_N[59] dyn2_dataIn_N[5] dyn2_dataIn_N[60] dyn2_dataIn_N[61] dyn2_dataIn_N[62]
+ dyn2_dataIn_N[63] dyn2_dataIn_N[6] dyn2_dataIn_N[7] dyn2_dataIn_N[8] dyn2_dataIn_N[9]
+ dyn2_dataIn_S[0] dyn2_dataIn_S[10] dyn2_dataIn_S[11] dyn2_dataIn_S[12] dyn2_dataIn_S[13]
+ dyn2_dataIn_S[14] dyn2_dataIn_S[15] dyn2_dataIn_S[16] dyn2_dataIn_S[17] dyn2_dataIn_S[18]
+ dyn2_dataIn_S[19] dyn2_dataIn_S[1] dyn2_dataIn_S[20] dyn2_dataIn_S[21] dyn2_dataIn_S[22]
+ dyn2_dataIn_S[23] dyn2_dataIn_S[24] dyn2_dataIn_S[25] dyn2_dataIn_S[26] dyn2_dataIn_S[27]
+ dyn2_dataIn_S[28] dyn2_dataIn_S[29] dyn2_dataIn_S[2] dyn2_dataIn_S[30] dyn2_dataIn_S[31]
+ dyn2_dataIn_S[32] dyn2_dataIn_S[33] dyn2_dataIn_S[34] dyn2_dataIn_S[35] dyn2_dataIn_S[36]
+ dyn2_dataIn_S[37] dyn2_dataIn_S[38] dyn2_dataIn_S[39] dyn2_dataIn_S[3] dyn2_dataIn_S[40]
+ dyn2_dataIn_S[41] dyn2_dataIn_S[42] dyn2_dataIn_S[43] dyn2_dataIn_S[44] dyn2_dataIn_S[45]
+ dyn2_dataIn_S[46] dyn2_dataIn_S[47] dyn2_dataIn_S[48] dyn2_dataIn_S[49] dyn2_dataIn_S[4]
+ dyn2_dataIn_S[50] dyn2_dataIn_S[51] dyn2_dataIn_S[52] dyn2_dataIn_S[53] dyn2_dataIn_S[54]
+ dyn2_dataIn_S[55] dyn2_dataIn_S[56] dyn2_dataIn_S[57] dyn2_dataIn_S[58] dyn2_dataIn_S[59]
+ dyn2_dataIn_S[5] dyn2_dataIn_S[60] dyn2_dataIn_S[61] dyn2_dataIn_S[62] dyn2_dataIn_S[63]
+ dyn2_dataIn_S[6] dyn2_dataIn_S[7] dyn2_dataIn_S[8] dyn2_dataIn_S[9] dyn2_dataIn_W[0]
+ dyn2_dataIn_W[10] dyn2_dataIn_W[11] dyn2_dataIn_W[12] dyn2_dataIn_W[13] dyn2_dataIn_W[14]
+ dyn2_dataIn_W[15] dyn2_dataIn_W[16] dyn2_dataIn_W[17] dyn2_dataIn_W[18] dyn2_dataIn_W[19]
+ dyn2_dataIn_W[1] dyn2_dataIn_W[20] dyn2_dataIn_W[21] dyn2_dataIn_W[22] dyn2_dataIn_W[23]
+ dyn2_dataIn_W[24] dyn2_dataIn_W[25] dyn2_dataIn_W[26] dyn2_dataIn_W[27] dyn2_dataIn_W[28]
+ dyn2_dataIn_W[29] dyn2_dataIn_W[2] dyn2_dataIn_W[30] dyn2_dataIn_W[31] dyn2_dataIn_W[32]
+ dyn2_dataIn_W[33] dyn2_dataIn_W[34] dyn2_dataIn_W[35] dyn2_dataIn_W[36] dyn2_dataIn_W[37]
+ dyn2_dataIn_W[38] dyn2_dataIn_W[39] dyn2_dataIn_W[3] dyn2_dataIn_W[40] dyn2_dataIn_W[41]
+ dyn2_dataIn_W[42] dyn2_dataIn_W[43] dyn2_dataIn_W[44] dyn2_dataIn_W[45] dyn2_dataIn_W[46]
+ dyn2_dataIn_W[47] dyn2_dataIn_W[48] dyn2_dataIn_W[49] dyn2_dataIn_W[4] dyn2_dataIn_W[50]
+ dyn2_dataIn_W[51] dyn2_dataIn_W[52] dyn2_dataIn_W[53] dyn2_dataIn_W[54] dyn2_dataIn_W[55]
+ dyn2_dataIn_W[56] dyn2_dataIn_W[57] dyn2_dataIn_W[58] dyn2_dataIn_W[59] dyn2_dataIn_W[5]
+ dyn2_dataIn_W[60] dyn2_dataIn_W[61] dyn2_dataIn_W[62] dyn2_dataIn_W[63] dyn2_dataIn_W[6]
+ dyn2_dataIn_W[7] dyn2_dataIn_W[8] dyn2_dataIn_W[9] dyn2_validIn_E dyn2_validIn_N
+ dyn2_validIn_S dyn2_validIn_W dyn2_yummyOut_E dyn2_yummyOut_N dyn2_yummyOut_S dyn2_yummyOut_W
+ flat_tileid[0] flat_tileid[1] flat_tileid[2] flat_tileid[3] flat_tileid[4] flat_tileid[5]
+ flat_tileid[6] flat_tileid[7] jtag_tiles_ucb_data[0] jtag_tiles_ucb_data[1] jtag_tiles_ucb_data[2]
+ jtag_tiles_ucb_data[3] jtag_tiles_ucb_val l15_config_req_address_s2[10] l15_config_req_address_s2[11]
+ l15_config_req_address_s2[12] l15_config_req_address_s2[13] l15_config_req_address_s2[14]
+ l15_config_req_address_s2[15] l15_config_req_address_s2[8] l15_config_req_address_s2[9]
+ l15_config_req_rw_s2 l15_config_req_val_s2 l15_config_write_req_data_s2[0] l15_config_write_req_data_s2[10]
+ l15_config_write_req_data_s2[11] l15_config_write_req_data_s2[12] l15_config_write_req_data_s2[13]
+ l15_config_write_req_data_s2[14] l15_config_write_req_data_s2[15] l15_config_write_req_data_s2[16]
+ l15_config_write_req_data_s2[17] l15_config_write_req_data_s2[18] l15_config_write_req_data_s2[19]
+ l15_config_write_req_data_s2[1] l15_config_write_req_data_s2[20] l15_config_write_req_data_s2[21]
+ l15_config_write_req_data_s2[22] l15_config_write_req_data_s2[23] l15_config_write_req_data_s2[24]
+ l15_config_write_req_data_s2[25] l15_config_write_req_data_s2[26] l15_config_write_req_data_s2[27]
+ l15_config_write_req_data_s2[28] l15_config_write_req_data_s2[29] l15_config_write_req_data_s2[2]
+ l15_config_write_req_data_s2[30] l15_config_write_req_data_s2[31] l15_config_write_req_data_s2[32]
+ l15_config_write_req_data_s2[33] l15_config_write_req_data_s2[34] l15_config_write_req_data_s2[35]
+ l15_config_write_req_data_s2[36] l15_config_write_req_data_s2[37] l15_config_write_req_data_s2[38]
+ l15_config_write_req_data_s2[39] l15_config_write_req_data_s2[3] l15_config_write_req_data_s2[40]
+ l15_config_write_req_data_s2[41] l15_config_write_req_data_s2[42] l15_config_write_req_data_s2[43]
+ l15_config_write_req_data_s2[44] l15_config_write_req_data_s2[45] l15_config_write_req_data_s2[46]
+ l15_config_write_req_data_s2[47] l15_config_write_req_data_s2[48] l15_config_write_req_data_s2[49]
+ l15_config_write_req_data_s2[4] l15_config_write_req_data_s2[50] l15_config_write_req_data_s2[51]
+ l15_config_write_req_data_s2[52] l15_config_write_req_data_s2[53] l15_config_write_req_data_s2[54]
+ l15_config_write_req_data_s2[55] l15_config_write_req_data_s2[56] l15_config_write_req_data_s2[57]
+ l15_config_write_req_data_s2[58] l15_config_write_req_data_s2[59] l15_config_write_req_data_s2[5]
+ l15_config_write_req_data_s2[60] l15_config_write_req_data_s2[61] l15_config_write_req_data_s2[62]
+ l15_config_write_req_data_s2[63] l15_config_write_req_data_s2[6] l15_config_write_req_data_s2[7]
+ l15_config_write_req_data_s2[8] l15_config_write_req_data_s2[9] l15_dmbr_l1missIn
+ l15_dmbr_l1missTag[0] l15_dmbr_l1missTag[1] l15_dmbr_l1missTag[2] l15_dmbr_l1missTag[3]
+ l15_dmbr_l2missIn l15_dmbr_l2missTag[0] l15_dmbr_l2missTag[1] l15_dmbr_l2missTag[2]
+ l15_dmbr_l2missTag[3] l15_dmbr_l2responseIn l15_transducer_ack l15_transducer_atomic
+ l15_transducer_blockinitstore l15_transducer_cross_invalidate l15_transducer_cross_invalidate_way[0]
+ l15_transducer_cross_invalidate_way[1] l15_transducer_data_0[0] l15_transducer_data_0[10]
+ l15_transducer_data_0[11] l15_transducer_data_0[12] l15_transducer_data_0[13] l15_transducer_data_0[14]
+ l15_transducer_data_0[15] l15_transducer_data_0[16] l15_transducer_data_0[17] l15_transducer_data_0[18]
+ l15_transducer_data_0[19] l15_transducer_data_0[1] l15_transducer_data_0[20] l15_transducer_data_0[21]
+ l15_transducer_data_0[22] l15_transducer_data_0[23] l15_transducer_data_0[24] l15_transducer_data_0[25]
+ l15_transducer_data_0[26] l15_transducer_data_0[27] l15_transducer_data_0[28] l15_transducer_data_0[29]
+ l15_transducer_data_0[2] l15_transducer_data_0[30] l15_transducer_data_0[31] l15_transducer_data_0[32]
+ l15_transducer_data_0[33] l15_transducer_data_0[34] l15_transducer_data_0[35] l15_transducer_data_0[36]
+ l15_transducer_data_0[37] l15_transducer_data_0[38] l15_transducer_data_0[39] l15_transducer_data_0[3]
+ l15_transducer_data_0[40] l15_transducer_data_0[41] l15_transducer_data_0[42] l15_transducer_data_0[43]
+ l15_transducer_data_0[44] l15_transducer_data_0[45] l15_transducer_data_0[46] l15_transducer_data_0[47]
+ l15_transducer_data_0[48] l15_transducer_data_0[49] l15_transducer_data_0[4] l15_transducer_data_0[50]
+ l15_transducer_data_0[51] l15_transducer_data_0[52] l15_transducer_data_0[53] l15_transducer_data_0[54]
+ l15_transducer_data_0[55] l15_transducer_data_0[56] l15_transducer_data_0[57] l15_transducer_data_0[58]
+ l15_transducer_data_0[59] l15_transducer_data_0[5] l15_transducer_data_0[60] l15_transducer_data_0[61]
+ l15_transducer_data_0[62] l15_transducer_data_0[63] l15_transducer_data_0[6] l15_transducer_data_0[7]
+ l15_transducer_data_0[8] l15_transducer_data_0[9] l15_transducer_data_1[0] l15_transducer_data_1[10]
+ l15_transducer_data_1[11] l15_transducer_data_1[12] l15_transducer_data_1[13] l15_transducer_data_1[14]
+ l15_transducer_data_1[15] l15_transducer_data_1[16] l15_transducer_data_1[17] l15_transducer_data_1[18]
+ l15_transducer_data_1[19] l15_transducer_data_1[1] l15_transducer_data_1[20] l15_transducer_data_1[21]
+ l15_transducer_data_1[22] l15_transducer_data_1[23] l15_transducer_data_1[24] l15_transducer_data_1[25]
+ l15_transducer_data_1[26] l15_transducer_data_1[27] l15_transducer_data_1[28] l15_transducer_data_1[29]
+ l15_transducer_data_1[2] l15_transducer_data_1[30] l15_transducer_data_1[31] l15_transducer_data_1[32]
+ l15_transducer_data_1[33] l15_transducer_data_1[34] l15_transducer_data_1[35] l15_transducer_data_1[36]
+ l15_transducer_data_1[37] l15_transducer_data_1[38] l15_transducer_data_1[39] l15_transducer_data_1[3]
+ l15_transducer_data_1[40] l15_transducer_data_1[41] l15_transducer_data_1[42] l15_transducer_data_1[43]
+ l15_transducer_data_1[44] l15_transducer_data_1[45] l15_transducer_data_1[46] l15_transducer_data_1[47]
+ l15_transducer_data_1[48] l15_transducer_data_1[49] l15_transducer_data_1[4] l15_transducer_data_1[50]
+ l15_transducer_data_1[51] l15_transducer_data_1[52] l15_transducer_data_1[53] l15_transducer_data_1[54]
+ l15_transducer_data_1[55] l15_transducer_data_1[56] l15_transducer_data_1[57] l15_transducer_data_1[58]
+ l15_transducer_data_1[59] l15_transducer_data_1[5] l15_transducer_data_1[60] l15_transducer_data_1[61]
+ l15_transducer_data_1[62] l15_transducer_data_1[63] l15_transducer_data_1[6] l15_transducer_data_1[7]
+ l15_transducer_data_1[8] l15_transducer_data_1[9] l15_transducer_data_2[0] l15_transducer_data_2[10]
+ l15_transducer_data_2[11] l15_transducer_data_2[12] l15_transducer_data_2[13] l15_transducer_data_2[14]
+ l15_transducer_data_2[15] l15_transducer_data_2[16] l15_transducer_data_2[17] l15_transducer_data_2[18]
+ l15_transducer_data_2[19] l15_transducer_data_2[1] l15_transducer_data_2[20] l15_transducer_data_2[21]
+ l15_transducer_data_2[22] l15_transducer_data_2[23] l15_transducer_data_2[24] l15_transducer_data_2[25]
+ l15_transducer_data_2[26] l15_transducer_data_2[27] l15_transducer_data_2[28] l15_transducer_data_2[29]
+ l15_transducer_data_2[2] l15_transducer_data_2[30] l15_transducer_data_2[31] l15_transducer_data_2[32]
+ l15_transducer_data_2[33] l15_transducer_data_2[34] l15_transducer_data_2[35] l15_transducer_data_2[36]
+ l15_transducer_data_2[37] l15_transducer_data_2[38] l15_transducer_data_2[39] l15_transducer_data_2[3]
+ l15_transducer_data_2[40] l15_transducer_data_2[41] l15_transducer_data_2[42] l15_transducer_data_2[43]
+ l15_transducer_data_2[44] l15_transducer_data_2[45] l15_transducer_data_2[46] l15_transducer_data_2[47]
+ l15_transducer_data_2[48] l15_transducer_data_2[49] l15_transducer_data_2[4] l15_transducer_data_2[50]
+ l15_transducer_data_2[51] l15_transducer_data_2[52] l15_transducer_data_2[53] l15_transducer_data_2[54]
+ l15_transducer_data_2[55] l15_transducer_data_2[56] l15_transducer_data_2[57] l15_transducer_data_2[58]
+ l15_transducer_data_2[59] l15_transducer_data_2[5] l15_transducer_data_2[60] l15_transducer_data_2[61]
+ l15_transducer_data_2[62] l15_transducer_data_2[63] l15_transducer_data_2[6] l15_transducer_data_2[7]
+ l15_transducer_data_2[8] l15_transducer_data_2[9] l15_transducer_data_3[0] l15_transducer_data_3[10]
+ l15_transducer_data_3[11] l15_transducer_data_3[12] l15_transducer_data_3[13] l15_transducer_data_3[14]
+ l15_transducer_data_3[15] l15_transducer_data_3[16] l15_transducer_data_3[17] l15_transducer_data_3[18]
+ l15_transducer_data_3[19] l15_transducer_data_3[1] l15_transducer_data_3[20] l15_transducer_data_3[21]
+ l15_transducer_data_3[22] l15_transducer_data_3[23] l15_transducer_data_3[24] l15_transducer_data_3[25]
+ l15_transducer_data_3[26] l15_transducer_data_3[27] l15_transducer_data_3[28] l15_transducer_data_3[29]
+ l15_transducer_data_3[2] l15_transducer_data_3[30] l15_transducer_data_3[31] l15_transducer_data_3[32]
+ l15_transducer_data_3[33] l15_transducer_data_3[34] l15_transducer_data_3[35] l15_transducer_data_3[36]
+ l15_transducer_data_3[37] l15_transducer_data_3[38] l15_transducer_data_3[39] l15_transducer_data_3[3]
+ l15_transducer_data_3[40] l15_transducer_data_3[41] l15_transducer_data_3[42] l15_transducer_data_3[43]
+ l15_transducer_data_3[44] l15_transducer_data_3[45] l15_transducer_data_3[46] l15_transducer_data_3[47]
+ l15_transducer_data_3[48] l15_transducer_data_3[49] l15_transducer_data_3[4] l15_transducer_data_3[50]
+ l15_transducer_data_3[51] l15_transducer_data_3[52] l15_transducer_data_3[53] l15_transducer_data_3[54]
+ l15_transducer_data_3[55] l15_transducer_data_3[56] l15_transducer_data_3[57] l15_transducer_data_3[58]
+ l15_transducer_data_3[59] l15_transducer_data_3[5] l15_transducer_data_3[60] l15_transducer_data_3[61]
+ l15_transducer_data_3[62] l15_transducer_data_3[63] l15_transducer_data_3[6] l15_transducer_data_3[7]
+ l15_transducer_data_3[8] l15_transducer_data_3[9] l15_transducer_error[0] l15_transducer_error[1]
+ l15_transducer_f4b l15_transducer_header_ack l15_transducer_inval_address_15_4[10]
+ l15_transducer_inval_address_15_4[11] l15_transducer_inval_address_15_4[12] l15_transducer_inval_address_15_4[13]
+ l15_transducer_inval_address_15_4[14] l15_transducer_inval_address_15_4[15] l15_transducer_inval_address_15_4[4]
+ l15_transducer_inval_address_15_4[5] l15_transducer_inval_address_15_4[6] l15_transducer_inval_address_15_4[7]
+ l15_transducer_inval_address_15_4[8] l15_transducer_inval_address_15_4[9] l15_transducer_inval_dcache_all_way
+ l15_transducer_inval_dcache_inval l15_transducer_inval_icache_all_way l15_transducer_inval_icache_inval
+ l15_transducer_inval_way[0] l15_transducer_inval_way[1] l15_transducer_l2miss l15_transducer_noncacheable
+ l15_transducer_prefetch l15_transducer_returntype[0] l15_transducer_returntype[1]
+ l15_transducer_returntype[2] l15_transducer_returntype[3] l15_transducer_threadid
+ l15_transducer_val l2_rtap_data[0] l2_rtap_data[1] l2_rtap_data[2] l2_rtap_data[3]
+ noc1_out_data[0] noc1_out_data[10] noc1_out_data[11] noc1_out_data[12] noc1_out_data[13]
+ noc1_out_data[14] noc1_out_data[15] noc1_out_data[16] noc1_out_data[17] noc1_out_data[18]
+ noc1_out_data[19] noc1_out_data[1] noc1_out_data[20] noc1_out_data[21] noc1_out_data[22]
+ noc1_out_data[23] noc1_out_data[24] noc1_out_data[25] noc1_out_data[26] noc1_out_data[27]
+ noc1_out_data[28] noc1_out_data[29] noc1_out_data[2] noc1_out_data[30] noc1_out_data[31]
+ noc1_out_data[32] noc1_out_data[33] noc1_out_data[34] noc1_out_data[35] noc1_out_data[36]
+ noc1_out_data[37] noc1_out_data[38] noc1_out_data[39] noc1_out_data[3] noc1_out_data[40]
+ noc1_out_data[41] noc1_out_data[42] noc1_out_data[43] noc1_out_data[44] noc1_out_data[45]
+ noc1_out_data[46] noc1_out_data[47] noc1_out_data[48] noc1_out_data[49] noc1_out_data[4]
+ noc1_out_data[50] noc1_out_data[51] noc1_out_data[52] noc1_out_data[53] noc1_out_data[54]
+ noc1_out_data[55] noc1_out_data[56] noc1_out_data[57] noc1_out_data[58] noc1_out_data[59]
+ noc1_out_data[5] noc1_out_data[60] noc1_out_data[61] noc1_out_data[62] noc1_out_data[63]
+ noc1_out_data[6] noc1_out_data[7] noc1_out_data[8] noc1_out_data[9] noc1_out_rdy
+ noc1_out_val noc2_in_data[0] noc2_in_data[10] noc2_in_data[11] noc2_in_data[12]
+ noc2_in_data[13] noc2_in_data[14] noc2_in_data[15] noc2_in_data[16] noc2_in_data[17]
+ noc2_in_data[18] noc2_in_data[19] noc2_in_data[1] noc2_in_data[20] noc2_in_data[21]
+ noc2_in_data[22] noc2_in_data[23] noc2_in_data[24] noc2_in_data[25] noc2_in_data[26]
+ noc2_in_data[27] noc2_in_data[28] noc2_in_data[29] noc2_in_data[2] noc2_in_data[30]
+ noc2_in_data[31] noc2_in_data[32] noc2_in_data[33] noc2_in_data[34] noc2_in_data[35]
+ noc2_in_data[36] noc2_in_data[37] noc2_in_data[38] noc2_in_data[39] noc2_in_data[3]
+ noc2_in_data[40] noc2_in_data[41] noc2_in_data[42] noc2_in_data[43] noc2_in_data[44]
+ noc2_in_data[45] noc2_in_data[46] noc2_in_data[47] noc2_in_data[48] noc2_in_data[49]
+ noc2_in_data[4] noc2_in_data[50] noc2_in_data[51] noc2_in_data[52] noc2_in_data[53]
+ noc2_in_data[54] noc2_in_data[55] noc2_in_data[56] noc2_in_data[57] noc2_in_data[58]
+ noc2_in_data[59] noc2_in_data[5] noc2_in_data[60] noc2_in_data[61] noc2_in_data[62]
+ noc2_in_data[63] noc2_in_data[6] noc2_in_data[7] noc2_in_data[8] noc2_in_data[9]
+ noc2_in_rdy noc2_in_val noc3_out_data[0] noc3_out_data[10] noc3_out_data[11] noc3_out_data[12]
+ noc3_out_data[13] noc3_out_data[14] noc3_out_data[15] noc3_out_data[16] noc3_out_data[17]
+ noc3_out_data[18] noc3_out_data[19] noc3_out_data[1] noc3_out_data[20] noc3_out_data[21]
+ noc3_out_data[22] noc3_out_data[23] noc3_out_data[24] noc3_out_data[25] noc3_out_data[26]
+ noc3_out_data[27] noc3_out_data[28] noc3_out_data[29] noc3_out_data[2] noc3_out_data[30]
+ noc3_out_data[31] noc3_out_data[32] noc3_out_data[33] noc3_out_data[34] noc3_out_data[35]
+ noc3_out_data[36] noc3_out_data[37] noc3_out_data[38] noc3_out_data[39] noc3_out_data[3]
+ noc3_out_data[40] noc3_out_data[41] noc3_out_data[42] noc3_out_data[43] noc3_out_data[44]
+ noc3_out_data[45] noc3_out_data[46] noc3_out_data[47] noc3_out_data[48] noc3_out_data[49]
+ noc3_out_data[4] noc3_out_data[50] noc3_out_data[51] noc3_out_data[52] noc3_out_data[53]
+ noc3_out_data[54] noc3_out_data[55] noc3_out_data[56] noc3_out_data[57] noc3_out_data[58]
+ noc3_out_data[59] noc3_out_data[5] noc3_out_data[60] noc3_out_data[61] noc3_out_data[62]
+ noc3_out_data[63] noc3_out_data[6] noc3_out_data[7] noc3_out_data[8] noc3_out_data[9]
+ noc3_out_rdy noc3_out_val processor_router_data_noc2[0] processor_router_data_noc2[10]
+ processor_router_data_noc2[11] processor_router_data_noc2[12] processor_router_data_noc2[13]
+ processor_router_data_noc2[14] processor_router_data_noc2[15] processor_router_data_noc2[16]
+ processor_router_data_noc2[17] processor_router_data_noc2[18] processor_router_data_noc2[19]
+ processor_router_data_noc2[1] processor_router_data_noc2[20] processor_router_data_noc2[21]
+ processor_router_data_noc2[22] processor_router_data_noc2[23] processor_router_data_noc2[24]
+ processor_router_data_noc2[25] processor_router_data_noc2[26] processor_router_data_noc2[27]
+ processor_router_data_noc2[28] processor_router_data_noc2[29] processor_router_data_noc2[2]
+ processor_router_data_noc2[30] processor_router_data_noc2[31] processor_router_data_noc2[32]
+ processor_router_data_noc2[33] processor_router_data_noc2[34] processor_router_data_noc2[35]
+ processor_router_data_noc2[36] processor_router_data_noc2[37] processor_router_data_noc2[38]
+ processor_router_data_noc2[39] processor_router_data_noc2[3] processor_router_data_noc2[40]
+ processor_router_data_noc2[41] processor_router_data_noc2[42] processor_router_data_noc2[43]
+ processor_router_data_noc2[44] processor_router_data_noc2[45] processor_router_data_noc2[46]
+ processor_router_data_noc2[47] processor_router_data_noc2[48] processor_router_data_noc2[49]
+ processor_router_data_noc2[4] processor_router_data_noc2[50] processor_router_data_noc2[51]
+ processor_router_data_noc2[52] processor_router_data_noc2[53] processor_router_data_noc2[54]
+ processor_router_data_noc2[55] processor_router_data_noc2[56] processor_router_data_noc2[57]
+ processor_router_data_noc2[58] processor_router_data_noc2[59] processor_router_data_noc2[5]
+ processor_router_data_noc2[60] processor_router_data_noc2[61] processor_router_data_noc2[62]
+ processor_router_data_noc2[63] processor_router_data_noc2[6] processor_router_data_noc2[7]
+ processor_router_data_noc2[8] processor_router_data_noc2[9] processor_router_ready_noc1
+ processor_router_ready_noc3 processor_router_valid_noc2 router_processor_ready_noc2
+ rst_n rtap_srams_bist_command[0] rtap_srams_bist_command[1] rtap_srams_bist_command[2]
+ rtap_srams_bist_command[3] rtap_srams_bist_data[0] rtap_srams_bist_data[1] rtap_srams_bist_data[2]
+ rtap_srams_bist_data[3] srams_rtap_data[0] srams_rtap_data[1] srams_rtap_data[2]
+ srams_rtap_data[3] tile_jtag_ucb_data[0] tile_jtag_ucb_data[1] tile_jtag_ucb_data[2]
+ tile_jtag_ucb_data[3] tile_jtag_ucb_val transducer_l15_address[0] transducer_l15_address[10]
+ transducer_l15_address[11] transducer_l15_address[12] transducer_l15_address[13]
+ transducer_l15_address[14] transducer_l15_address[15] transducer_l15_address[16]
+ transducer_l15_address[17] transducer_l15_address[18] transducer_l15_address[19]
+ transducer_l15_address[1] transducer_l15_address[20] transducer_l15_address[21]
+ transducer_l15_address[22] transducer_l15_address[23] transducer_l15_address[24]
+ transducer_l15_address[25] transducer_l15_address[26] transducer_l15_address[27]
+ transducer_l15_address[28] transducer_l15_address[29] transducer_l15_address[2]
+ transducer_l15_address[30] transducer_l15_address[31] transducer_l15_address[32]
+ transducer_l15_address[33] transducer_l15_address[34] transducer_l15_address[35]
+ transducer_l15_address[36] transducer_l15_address[37] transducer_l15_address[38]
+ transducer_l15_address[39] transducer_l15_address[3] transducer_l15_address[4] transducer_l15_address[5]
+ transducer_l15_address[6] transducer_l15_address[7] transducer_l15_address[8] transducer_l15_address[9]
+ transducer_l15_amo_op[0] transducer_l15_amo_op[1] transducer_l15_amo_op[2] transducer_l15_amo_op[3]
+ transducer_l15_blockinitstore transducer_l15_blockstore transducer_l15_csm_data[0]
+ transducer_l15_csm_data[10] transducer_l15_csm_data[11] transducer_l15_csm_data[12]
+ transducer_l15_csm_data[13] transducer_l15_csm_data[14] transducer_l15_csm_data[15]
+ transducer_l15_csm_data[16] transducer_l15_csm_data[17] transducer_l15_csm_data[18]
+ transducer_l15_csm_data[19] transducer_l15_csm_data[1] transducer_l15_csm_data[20]
+ transducer_l15_csm_data[21] transducer_l15_csm_data[22] transducer_l15_csm_data[23]
+ transducer_l15_csm_data[24] transducer_l15_csm_data[25] transducer_l15_csm_data[26]
+ transducer_l15_csm_data[27] transducer_l15_csm_data[28] transducer_l15_csm_data[29]
+ transducer_l15_csm_data[2] transducer_l15_csm_data[30] transducer_l15_csm_data[31]
+ transducer_l15_csm_data[32] transducer_l15_csm_data[3] transducer_l15_csm_data[4]
+ transducer_l15_csm_data[5] transducer_l15_csm_data[6] transducer_l15_csm_data[7]
+ transducer_l15_csm_data[8] transducer_l15_csm_data[9] transducer_l15_data[0] transducer_l15_data[10]
+ transducer_l15_data[11] transducer_l15_data[12] transducer_l15_data[13] transducer_l15_data[14]
+ transducer_l15_data[15] transducer_l15_data[16] transducer_l15_data[17] transducer_l15_data[18]
+ transducer_l15_data[19] transducer_l15_data[1] transducer_l15_data[20] transducer_l15_data[21]
+ transducer_l15_data[22] transducer_l15_data[23] transducer_l15_data[24] transducer_l15_data[25]
+ transducer_l15_data[26] transducer_l15_data[27] transducer_l15_data[28] transducer_l15_data[29]
+ transducer_l15_data[2] transducer_l15_data[30] transducer_l15_data[31] transducer_l15_data[32]
+ transducer_l15_data[33] transducer_l15_data[34] transducer_l15_data[35] transducer_l15_data[36]
+ transducer_l15_data[37] transducer_l15_data[38] transducer_l15_data[39] transducer_l15_data[3]
+ transducer_l15_data[40] transducer_l15_data[41] transducer_l15_data[42] transducer_l15_data[43]
+ transducer_l15_data[44] transducer_l15_data[45] transducer_l15_data[46] transducer_l15_data[47]
+ transducer_l15_data[48] transducer_l15_data[49] transducer_l15_data[4] transducer_l15_data[50]
+ transducer_l15_data[51] transducer_l15_data[52] transducer_l15_data[53] transducer_l15_data[54]
+ transducer_l15_data[55] transducer_l15_data[56] transducer_l15_data[57] transducer_l15_data[58]
+ transducer_l15_data[59] transducer_l15_data[5] transducer_l15_data[60] transducer_l15_data[61]
+ transducer_l15_data[62] transducer_l15_data[63] transducer_l15_data[6] transducer_l15_data[7]
+ transducer_l15_data[8] transducer_l15_data[9] transducer_l15_data_next_entry[0]
+ transducer_l15_data_next_entry[10] transducer_l15_data_next_entry[11] transducer_l15_data_next_entry[12]
+ transducer_l15_data_next_entry[13] transducer_l15_data_next_entry[14] transducer_l15_data_next_entry[15]
+ transducer_l15_data_next_entry[16] transducer_l15_data_next_entry[17] transducer_l15_data_next_entry[18]
+ transducer_l15_data_next_entry[19] transducer_l15_data_next_entry[1] transducer_l15_data_next_entry[20]
+ transducer_l15_data_next_entry[21] transducer_l15_data_next_entry[22] transducer_l15_data_next_entry[23]
+ transducer_l15_data_next_entry[24] transducer_l15_data_next_entry[25] transducer_l15_data_next_entry[26]
+ transducer_l15_data_next_entry[27] transducer_l15_data_next_entry[28] transducer_l15_data_next_entry[29]
+ transducer_l15_data_next_entry[2] transducer_l15_data_next_entry[30] transducer_l15_data_next_entry[31]
+ transducer_l15_data_next_entry[32] transducer_l15_data_next_entry[33] transducer_l15_data_next_entry[34]
+ transducer_l15_data_next_entry[35] transducer_l15_data_next_entry[36] transducer_l15_data_next_entry[37]
+ transducer_l15_data_next_entry[38] transducer_l15_data_next_entry[39] transducer_l15_data_next_entry[3]
+ transducer_l15_data_next_entry[40] transducer_l15_data_next_entry[41] transducer_l15_data_next_entry[42]
+ transducer_l15_data_next_entry[43] transducer_l15_data_next_entry[44] transducer_l15_data_next_entry[45]
+ transducer_l15_data_next_entry[46] transducer_l15_data_next_entry[47] transducer_l15_data_next_entry[48]
+ transducer_l15_data_next_entry[49] transducer_l15_data_next_entry[4] transducer_l15_data_next_entry[50]
+ transducer_l15_data_next_entry[51] transducer_l15_data_next_entry[52] transducer_l15_data_next_entry[53]
+ transducer_l15_data_next_entry[54] transducer_l15_data_next_entry[55] transducer_l15_data_next_entry[56]
+ transducer_l15_data_next_entry[57] transducer_l15_data_next_entry[58] transducer_l15_data_next_entry[59]
+ transducer_l15_data_next_entry[5] transducer_l15_data_next_entry[60] transducer_l15_data_next_entry[61]
+ transducer_l15_data_next_entry[62] transducer_l15_data_next_entry[63] transducer_l15_data_next_entry[6]
+ transducer_l15_data_next_entry[7] transducer_l15_data_next_entry[8] transducer_l15_data_next_entry[9]
+ transducer_l15_invalidate_cacheline transducer_l15_l1rplway[0] transducer_l15_l1rplway[1]
+ transducer_l15_nc transducer_l15_prefetch transducer_l15_req_ack transducer_l15_rqtype[0]
+ transducer_l15_rqtype[1] transducer_l15_rqtype[2] transducer_l15_rqtype[3] transducer_l15_rqtype[4]
+ transducer_l15_size[0] transducer_l15_size[1] transducer_l15_size[2] transducer_l15_threadid
+ transducer_l15_val vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xtile tile/buffer_processor_data_noc1[0] tile/buffer_processor_data_noc1[10] tile/buffer_processor_data_noc1[11]
+ tile/buffer_processor_data_noc1[12] tile/buffer_processor_data_noc1[13] tile/buffer_processor_data_noc1[14]
+ tile/buffer_processor_data_noc1[15] tile/buffer_processor_data_noc1[16] tile/buffer_processor_data_noc1[17]
+ tile/buffer_processor_data_noc1[18] tile/buffer_processor_data_noc1[19] tile/buffer_processor_data_noc1[1]
+ tile/buffer_processor_data_noc1[20] tile/buffer_processor_data_noc1[21] tile/buffer_processor_data_noc1[22]
+ tile/buffer_processor_data_noc1[23] tile/buffer_processor_data_noc1[24] tile/buffer_processor_data_noc1[25]
+ tile/buffer_processor_data_noc1[26] tile/buffer_processor_data_noc1[27] tile/buffer_processor_data_noc1[28]
+ tile/buffer_processor_data_noc1[29] tile/buffer_processor_data_noc1[2] tile/buffer_processor_data_noc1[30]
+ tile/buffer_processor_data_noc1[31] tile/buffer_processor_data_noc1[32] tile/buffer_processor_data_noc1[33]
+ tile/buffer_processor_data_noc1[34] tile/buffer_processor_data_noc1[35] tile/buffer_processor_data_noc1[36]
+ tile/buffer_processor_data_noc1[37] tile/buffer_processor_data_noc1[38] tile/buffer_processor_data_noc1[39]
+ tile/buffer_processor_data_noc1[3] tile/buffer_processor_data_noc1[40] tile/buffer_processor_data_noc1[41]
+ tile/buffer_processor_data_noc1[42] tile/buffer_processor_data_noc1[43] tile/buffer_processor_data_noc1[44]
+ tile/buffer_processor_data_noc1[45] tile/buffer_processor_data_noc1[46] tile/buffer_processor_data_noc1[47]
+ tile/buffer_processor_data_noc1[48] tile/buffer_processor_data_noc1[49] tile/buffer_processor_data_noc1[4]
+ tile/buffer_processor_data_noc1[50] tile/buffer_processor_data_noc1[51] tile/buffer_processor_data_noc1[52]
+ tile/buffer_processor_data_noc1[53] tile/buffer_processor_data_noc1[54] tile/buffer_processor_data_noc1[55]
+ tile/buffer_processor_data_noc1[56] tile/buffer_processor_data_noc1[57] tile/buffer_processor_data_noc1[58]
+ tile/buffer_processor_data_noc1[59] tile/buffer_processor_data_noc1[5] tile/buffer_processor_data_noc1[60]
+ tile/buffer_processor_data_noc1[61] tile/buffer_processor_data_noc1[62] tile/buffer_processor_data_noc1[63]
+ tile/buffer_processor_data_noc1[6] tile/buffer_processor_data_noc1[7] tile/buffer_processor_data_noc1[8]
+ tile/buffer_processor_data_noc1[9] tile/buffer_processor_data_noc3[0] tile/buffer_processor_data_noc3[10]
+ tile/buffer_processor_data_noc3[11] tile/buffer_processor_data_noc3[12] tile/buffer_processor_data_noc3[13]
+ tile/buffer_processor_data_noc3[14] tile/buffer_processor_data_noc3[15] tile/buffer_processor_data_noc3[16]
+ tile/buffer_processor_data_noc3[17] tile/buffer_processor_data_noc3[18] tile/buffer_processor_data_noc3[19]
+ tile/buffer_processor_data_noc3[1] tile/buffer_processor_data_noc3[20] tile/buffer_processor_data_noc3[21]
+ tile/buffer_processor_data_noc3[22] tile/buffer_processor_data_noc3[23] tile/buffer_processor_data_noc3[24]
+ tile/buffer_processor_data_noc3[25] tile/buffer_processor_data_noc3[26] tile/buffer_processor_data_noc3[27]
+ tile/buffer_processor_data_noc3[28] tile/buffer_processor_data_noc3[29] tile/buffer_processor_data_noc3[2]
+ tile/buffer_processor_data_noc3[30] tile/buffer_processor_data_noc3[31] tile/buffer_processor_data_noc3[32]
+ tile/buffer_processor_data_noc3[33] tile/buffer_processor_data_noc3[34] tile/buffer_processor_data_noc3[35]
+ tile/buffer_processor_data_noc3[36] tile/buffer_processor_data_noc3[37] tile/buffer_processor_data_noc3[38]
+ tile/buffer_processor_data_noc3[39] tile/buffer_processor_data_noc3[3] tile/buffer_processor_data_noc3[40]
+ tile/buffer_processor_data_noc3[41] tile/buffer_processor_data_noc3[42] tile/buffer_processor_data_noc3[43]
+ tile/buffer_processor_data_noc3[44] tile/buffer_processor_data_noc3[45] tile/buffer_processor_data_noc3[46]
+ tile/buffer_processor_data_noc3[47] tile/buffer_processor_data_noc3[48] tile/buffer_processor_data_noc3[49]
+ tile/buffer_processor_data_noc3[4] tile/buffer_processor_data_noc3[50] tile/buffer_processor_data_noc3[51]
+ tile/buffer_processor_data_noc3[52] tile/buffer_processor_data_noc3[53] tile/buffer_processor_data_noc3[54]
+ tile/buffer_processor_data_noc3[55] tile/buffer_processor_data_noc3[56] tile/buffer_processor_data_noc3[57]
+ tile/buffer_processor_data_noc3[58] tile/buffer_processor_data_noc3[59] tile/buffer_processor_data_noc3[5]
+ tile/buffer_processor_data_noc3[60] tile/buffer_processor_data_noc3[61] tile/buffer_processor_data_noc3[62]
+ tile/buffer_processor_data_noc3[63] tile/buffer_processor_data_noc3[6] tile/buffer_processor_data_noc3[7]
+ tile/buffer_processor_data_noc3[8] tile/buffer_processor_data_noc3[9] tile/buffer_processor_valid_noc1
+ tile/buffer_processor_valid_noc3 tile/chipid[0] tile/chipid[10] tile/chipid[11]
+ tile/chipid[12] tile/chipid[13] tile/chipid[1] tile/chipid[2] tile/chipid[3] tile/chipid[4]
+ tile/chipid[5] tile/chipid[6] tile/chipid[7] tile/chipid[8] tile/chipid[9] wb_clk_i
+ tile/clk_en tile/config_chipid[0] tile/config_chipid[10] tile/config_chipid[11]
+ tile/config_chipid[12] tile/config_chipid[13] tile/config_chipid[1] tile/config_chipid[2]
+ tile/config_chipid[3] tile/config_chipid[4] tile/config_chipid[5] tile/config_chipid[6]
+ tile/config_chipid[7] tile/config_chipid[8] tile/config_chipid[9] tile/config_coreid_x[0]
+ tile/config_coreid_x[1] tile/config_coreid_x[2] tile/config_coreid_x[3] tile/config_coreid_x[4]
+ tile/config_coreid_x[5] tile/config_coreid_x[6] tile/config_coreid_x[7] tile/config_coreid_y[0]
+ tile/config_coreid_y[1] tile/config_coreid_y[2] tile/config_coreid_y[3] tile/config_coreid_y[4]
+ tile/config_coreid_y[5] tile/config_coreid_y[6] tile/config_coreid_y[7] tile/config_csm_en
+ tile/config_hmt_base[0] tile/config_hmt_base[10] tile/config_hmt_base[11] tile/config_hmt_base[12]
+ tile/config_hmt_base[13] tile/config_hmt_base[14] tile/config_hmt_base[15] tile/config_hmt_base[16]
+ tile/config_hmt_base[17] tile/config_hmt_base[18] tile/config_hmt_base[19] tile/config_hmt_base[1]
+ tile/config_hmt_base[20] tile/config_hmt_base[21] tile/config_hmt_base[2] tile/config_hmt_base[3]
+ tile/config_hmt_base[4] tile/config_hmt_base[5] tile/config_hmt_base[6] tile/config_hmt_base[7]
+ tile/config_hmt_base[8] tile/config_hmt_base[9] tile/config_home_alloc_method[0]
+ tile/config_home_alloc_method[1] tile/config_l15_read_res_data_s3[0] tile/config_l15_read_res_data_s3[10]
+ tile/config_l15_read_res_data_s3[11] tile/config_l15_read_res_data_s3[12] tile/config_l15_read_res_data_s3[13]
+ tile/config_l15_read_res_data_s3[14] tile/config_l15_read_res_data_s3[15] tile/config_l15_read_res_data_s3[16]
+ tile/config_l15_read_res_data_s3[17] tile/config_l15_read_res_data_s3[18] tile/config_l15_read_res_data_s3[19]
+ tile/config_l15_read_res_data_s3[1] tile/config_l15_read_res_data_s3[20] tile/config_l15_read_res_data_s3[21]
+ tile/config_l15_read_res_data_s3[22] tile/config_l15_read_res_data_s3[23] tile/config_l15_read_res_data_s3[24]
+ tile/config_l15_read_res_data_s3[25] tile/config_l15_read_res_data_s3[26] tile/config_l15_read_res_data_s3[27]
+ tile/config_l15_read_res_data_s3[28] tile/config_l15_read_res_data_s3[29] tile/config_l15_read_res_data_s3[2]
+ tile/config_l15_read_res_data_s3[30] tile/config_l15_read_res_data_s3[31] tile/config_l15_read_res_data_s3[32]
+ tile/config_l15_read_res_data_s3[33] tile/config_l15_read_res_data_s3[34] tile/config_l15_read_res_data_s3[35]
+ tile/config_l15_read_res_data_s3[36] tile/config_l15_read_res_data_s3[37] tile/config_l15_read_res_data_s3[38]
+ tile/config_l15_read_res_data_s3[39] tile/config_l15_read_res_data_s3[3] tile/config_l15_read_res_data_s3[40]
+ tile/config_l15_read_res_data_s3[41] tile/config_l15_read_res_data_s3[42] tile/config_l15_read_res_data_s3[43]
+ tile/config_l15_read_res_data_s3[44] tile/config_l15_read_res_data_s3[45] tile/config_l15_read_res_data_s3[46]
+ tile/config_l15_read_res_data_s3[47] tile/config_l15_read_res_data_s3[48] tile/config_l15_read_res_data_s3[49]
+ tile/config_l15_read_res_data_s3[4] tile/config_l15_read_res_data_s3[50] tile/config_l15_read_res_data_s3[51]
+ tile/config_l15_read_res_data_s3[52] tile/config_l15_read_res_data_s3[53] tile/config_l15_read_res_data_s3[54]
+ tile/config_l15_read_res_data_s3[55] tile/config_l15_read_res_data_s3[56] tile/config_l15_read_res_data_s3[57]
+ tile/config_l15_read_res_data_s3[58] tile/config_l15_read_res_data_s3[59] tile/config_l15_read_res_data_s3[5]
+ tile/config_l15_read_res_data_s3[60] tile/config_l15_read_res_data_s3[61] tile/config_l15_read_res_data_s3[62]
+ tile/config_l15_read_res_data_s3[63] tile/config_l15_read_res_data_s3[6] tile/config_l15_read_res_data_s3[7]
+ tile/config_l15_read_res_data_s3[8] tile/config_l15_read_res_data_s3[9] tile/config_system_tile_count_5_0[0]
+ tile/config_system_tile_count_5_0[1] tile/config_system_tile_count_5_0[2] tile/config_system_tile_count_5_0[3]
+ tile/config_system_tile_count_5_0[4] tile/config_system_tile_count_5_0[5] tile/coreid_x[0]
+ tile/coreid_x[1] tile/coreid_x[2] tile/coreid_x[3] tile/coreid_x[4] tile/coreid_x[5]
+ tile/coreid_x[6] tile/coreid_x[7] tile/coreid_y[0] tile/coreid_y[1] tile/coreid_y[2]
+ tile/coreid_y[3] tile/coreid_y[4] tile/coreid_y[5] tile/coreid_y[6] tile/coreid_y[7]
+ tile/default_chipid[0] tile/default_chipid[10] tile/default_chipid[11] tile/default_chipid[12]
+ tile/default_chipid[13] tile/default_chipid[1] tile/default_chipid[2] tile/default_chipid[3]
+ tile/default_chipid[4] tile/default_chipid[5] tile/default_chipid[6] tile/default_chipid[7]
+ tile/default_chipid[8] tile/default_chipid[9] tile/default_coreid_x[0] tile/default_coreid_x[1]
+ tile/default_coreid_x[2] tile/default_coreid_x[3] tile/default_coreid_x[4] tile/default_coreid_x[5]
+ tile/default_coreid_x[6] tile/default_coreid_x[7] tile/default_coreid_y[0] tile/default_coreid_y[1]
+ tile/default_coreid_y[2] tile/default_coreid_y[3] tile/default_coreid_y[4] tile/default_coreid_y[5]
+ tile/default_coreid_y[6] tile/default_coreid_y[7] tile/dmbr_l15_stall tile/dummy_core[0]
+ tile/dummy_core[10] tile/dummy_core[11] tile/dummy_core[12] tile/dummy_core[13]
+ tile/dummy_core[14] tile/dummy_core[15] tile/dummy_core[16] tile/dummy_core[17]
+ tile/dummy_core[18] tile/dummy_core[19] tile/dummy_core[1] tile/dummy_core[20] tile/dummy_core[21]
+ tile/dummy_core[22] tile/dummy_core[23] tile/dummy_core[24] tile/dummy_core[25]
+ tile/dummy_core[26] tile/dummy_core[27] tile/dummy_core[28] tile/dummy_core[29]
+ tile/dummy_core[2] tile/dummy_core[30] tile/dummy_core[31] tile/dummy_core[3] tile/dummy_core[4]
+ tile/dummy_core[5] tile/dummy_core[6] tile/dummy_core[7] tile/dummy_core[8] tile/dummy_core[9]
+ tile/dyn0_dEo[0] tile/dyn0_dEo[10] tile/dyn0_dEo[11] tile/dyn0_dEo[12] tile/dyn0_dEo[13]
+ tile/dyn0_dEo[14] tile/dyn0_dEo[15] tile/dyn0_dEo[16] tile/dyn0_dEo[17] tile/dyn0_dEo[18]
+ tile/dyn0_dEo[19] tile/dyn0_dEo[1] tile/dyn0_dEo[20] tile/dyn0_dEo[21] tile/dyn0_dEo[22]
+ tile/dyn0_dEo[23] tile/dyn0_dEo[24] tile/dyn0_dEo[25] tile/dyn0_dEo[26] tile/dyn0_dEo[27]
+ tile/dyn0_dEo[28] tile/dyn0_dEo[29] tile/dyn0_dEo[2] tile/dyn0_dEo[30] tile/dyn0_dEo[31]
+ tile/dyn0_dEo[32] tile/dyn0_dEo[33] tile/dyn0_dEo[34] tile/dyn0_dEo[35] tile/dyn0_dEo[36]
+ tile/dyn0_dEo[37] tile/dyn0_dEo[38] tile/dyn0_dEo[39] tile/dyn0_dEo[3] tile/dyn0_dEo[40]
+ tile/dyn0_dEo[41] tile/dyn0_dEo[42] tile/dyn0_dEo[43] tile/dyn0_dEo[44] tile/dyn0_dEo[45]
+ tile/dyn0_dEo[46] tile/dyn0_dEo[47] tile/dyn0_dEo[48] tile/dyn0_dEo[49] tile/dyn0_dEo[4]
+ tile/dyn0_dEo[50] tile/dyn0_dEo[51] tile/dyn0_dEo[52] tile/dyn0_dEo[53] tile/dyn0_dEo[54]
+ tile/dyn0_dEo[55] tile/dyn0_dEo[56] tile/dyn0_dEo[57] tile/dyn0_dEo[58] tile/dyn0_dEo[59]
+ tile/dyn0_dEo[5] tile/dyn0_dEo[60] tile/dyn0_dEo[61] tile/dyn0_dEo[62] tile/dyn0_dEo[63]
+ tile/dyn0_dEo[6] tile/dyn0_dEo[7] tile/dyn0_dEo[8] tile/dyn0_dEo[9] io_out[1] tile/dyn0_dEo_yummy
+ tile/dyn0_dNo[0] tile/dyn0_dNo[10] tile/dyn0_dNo[11] tile/dyn0_dNo[12] tile/dyn0_dNo[13]
+ tile/dyn0_dNo[14] tile/dyn0_dNo[15] tile/dyn0_dNo[16] tile/dyn0_dNo[17] tile/dyn0_dNo[18]
+ tile/dyn0_dNo[19] tile/dyn0_dNo[1] tile/dyn0_dNo[20] tile/dyn0_dNo[21] tile/dyn0_dNo[22]
+ tile/dyn0_dNo[23] tile/dyn0_dNo[24] tile/dyn0_dNo[25] tile/dyn0_dNo[26] tile/dyn0_dNo[27]
+ tile/dyn0_dNo[28] tile/dyn0_dNo[29] tile/dyn0_dNo[2] tile/dyn0_dNo[30] tile/dyn0_dNo[31]
+ tile/dyn0_dNo[32] tile/dyn0_dNo[33] tile/dyn0_dNo[34] tile/dyn0_dNo[35] tile/dyn0_dNo[36]
+ tile/dyn0_dNo[37] tile/dyn0_dNo[38] tile/dyn0_dNo[39] tile/dyn0_dNo[3] tile/dyn0_dNo[40]
+ tile/dyn0_dNo[41] tile/dyn0_dNo[42] tile/dyn0_dNo[43] tile/dyn0_dNo[44] tile/dyn0_dNo[45]
+ tile/dyn0_dNo[46] tile/dyn0_dNo[47] tile/dyn0_dNo[48] tile/dyn0_dNo[49] tile/dyn0_dNo[4]
+ tile/dyn0_dNo[50] tile/dyn0_dNo[51] tile/dyn0_dNo[52] tile/dyn0_dNo[53] tile/dyn0_dNo[54]
+ tile/dyn0_dNo[55] tile/dyn0_dNo[56] tile/dyn0_dNo[57] tile/dyn0_dNo[58] tile/dyn0_dNo[59]
+ tile/dyn0_dNo[5] tile/dyn0_dNo[60] tile/dyn0_dNo[61] tile/dyn0_dNo[62] tile/dyn0_dNo[63]
+ tile/dyn0_dNo[6] tile/dyn0_dNo[7] tile/dyn0_dNo[8] tile/dyn0_dNo[9] io_out[0] tile/dyn0_dNo_yummy
+ tile/dyn0_dSo[0] tile/dyn0_dSo[10] tile/dyn0_dSo[11] tile/dyn0_dSo[12] tile/dyn0_dSo[13]
+ tile/dyn0_dSo[14] tile/dyn0_dSo[15] tile/dyn0_dSo[16] tile/dyn0_dSo[17] tile/dyn0_dSo[18]
+ tile/dyn0_dSo[19] tile/dyn0_dSo[1] tile/dyn0_dSo[20] tile/dyn0_dSo[21] tile/dyn0_dSo[22]
+ tile/dyn0_dSo[23] tile/dyn0_dSo[24] tile/dyn0_dSo[25] tile/dyn0_dSo[26] tile/dyn0_dSo[27]
+ tile/dyn0_dSo[28] tile/dyn0_dSo[29] tile/dyn0_dSo[2] tile/dyn0_dSo[30] tile/dyn0_dSo[31]
+ tile/dyn0_dSo[32] tile/dyn0_dSo[33] tile/dyn0_dSo[34] tile/dyn0_dSo[35] tile/dyn0_dSo[36]
+ tile/dyn0_dSo[37] tile/dyn0_dSo[38] tile/dyn0_dSo[39] tile/dyn0_dSo[3] tile/dyn0_dSo[40]
+ tile/dyn0_dSo[41] tile/dyn0_dSo[42] tile/dyn0_dSo[43] tile/dyn0_dSo[44] tile/dyn0_dSo[45]
+ tile/dyn0_dSo[46] tile/dyn0_dSo[47] tile/dyn0_dSo[48] tile/dyn0_dSo[49] tile/dyn0_dSo[4]
+ tile/dyn0_dSo[50] tile/dyn0_dSo[51] tile/dyn0_dSo[52] tile/dyn0_dSo[53] tile/dyn0_dSo[54]
+ tile/dyn0_dSo[55] tile/dyn0_dSo[56] tile/dyn0_dSo[57] tile/dyn0_dSo[58] tile/dyn0_dSo[59]
+ tile/dyn0_dSo[5] tile/dyn0_dSo[60] tile/dyn0_dSo[61] tile/dyn0_dSo[62] tile/dyn0_dSo[63]
+ tile/dyn0_dSo[6] tile/dyn0_dSo[7] tile/dyn0_dSo[8] tile/dyn0_dSo[9] io_out[3] tile/dyn0_dSo_yummy
+ tile/dyn0_dWo[0] tile/dyn0_dWo[10] tile/dyn0_dWo[11] tile/dyn0_dWo[12] tile/dyn0_dWo[13]
+ tile/dyn0_dWo[14] tile/dyn0_dWo[15] tile/dyn0_dWo[16] tile/dyn0_dWo[17] tile/dyn0_dWo[18]
+ tile/dyn0_dWo[19] tile/dyn0_dWo[1] tile/dyn0_dWo[20] tile/dyn0_dWo[21] tile/dyn0_dWo[22]
+ tile/dyn0_dWo[23] tile/dyn0_dWo[24] tile/dyn0_dWo[25] tile/dyn0_dWo[26] tile/dyn0_dWo[27]
+ tile/dyn0_dWo[28] tile/dyn0_dWo[29] tile/dyn0_dWo[2] tile/dyn0_dWo[30] tile/dyn0_dWo[31]
+ tile/dyn0_dWo[32] tile/dyn0_dWo[33] tile/dyn0_dWo[34] tile/dyn0_dWo[35] tile/dyn0_dWo[36]
+ tile/dyn0_dWo[37] tile/dyn0_dWo[38] tile/dyn0_dWo[39] tile/dyn0_dWo[3] tile/dyn0_dWo[40]
+ tile/dyn0_dWo[41] tile/dyn0_dWo[42] tile/dyn0_dWo[43] tile/dyn0_dWo[44] tile/dyn0_dWo[45]
+ tile/dyn0_dWo[46] tile/dyn0_dWo[47] tile/dyn0_dWo[48] tile/dyn0_dWo[49] tile/dyn0_dWo[4]
+ tile/dyn0_dWo[50] tile/dyn0_dWo[51] tile/dyn0_dWo[52] tile/dyn0_dWo[53] tile/dyn0_dWo[54]
+ tile/dyn0_dWo[55] tile/dyn0_dWo[56] tile/dyn0_dWo[57] tile/dyn0_dWo[58] tile/dyn0_dWo[59]
+ tile/dyn0_dWo[5] tile/dyn0_dWo[60] tile/dyn0_dWo[61] tile/dyn0_dWo[62] tile/dyn0_dWo[63]
+ tile/dyn0_dWo[6] tile/dyn0_dWo[7] tile/dyn0_dWo[8] tile/dyn0_dWo[9] io_out[2] tile/dyn0_dWo_yummy
+ tile/dyn0_dataIn_E[0] tile/dyn0_dataIn_E[10] tile/dyn0_dataIn_E[11] tile/dyn0_dataIn_E[12]
+ tile/dyn0_dataIn_E[13] tile/dyn0_dataIn_E[14] tile/dyn0_dataIn_E[15] tile/dyn0_dataIn_E[16]
+ tile/dyn0_dataIn_E[17] tile/dyn0_dataIn_E[18] tile/dyn0_dataIn_E[19] tile/dyn0_dataIn_E[1]
+ tile/dyn0_dataIn_E[20] tile/dyn0_dataIn_E[21] tile/dyn0_dataIn_E[22] tile/dyn0_dataIn_E[23]
+ tile/dyn0_dataIn_E[24] tile/dyn0_dataIn_E[25] tile/dyn0_dataIn_E[26] tile/dyn0_dataIn_E[27]
+ tile/dyn0_dataIn_E[28] tile/dyn0_dataIn_E[29] tile/dyn0_dataIn_E[2] tile/dyn0_dataIn_E[30]
+ tile/dyn0_dataIn_E[31] tile/dyn0_dataIn_E[32] tile/dyn0_dataIn_E[33] tile/dyn0_dataIn_E[34]
+ tile/dyn0_dataIn_E[35] tile/dyn0_dataIn_E[36] tile/dyn0_dataIn_E[37] tile/dyn0_dataIn_E[38]
+ tile/dyn0_dataIn_E[39] tile/dyn0_dataIn_E[3] tile/dyn0_dataIn_E[40] tile/dyn0_dataIn_E[41]
+ tile/dyn0_dataIn_E[42] tile/dyn0_dataIn_E[43] tile/dyn0_dataIn_E[44] tile/dyn0_dataIn_E[45]
+ tile/dyn0_dataIn_E[46] tile/dyn0_dataIn_E[47] tile/dyn0_dataIn_E[48] tile/dyn0_dataIn_E[49]
+ tile/dyn0_dataIn_E[4] tile/dyn0_dataIn_E[50] tile/dyn0_dataIn_E[51] tile/dyn0_dataIn_E[52]
+ tile/dyn0_dataIn_E[53] tile/dyn0_dataIn_E[54] tile/dyn0_dataIn_E[55] tile/dyn0_dataIn_E[56]
+ tile/dyn0_dataIn_E[57] tile/dyn0_dataIn_E[58] tile/dyn0_dataIn_E[59] tile/dyn0_dataIn_E[5]
+ tile/dyn0_dataIn_E[60] tile/dyn0_dataIn_E[61] tile/dyn0_dataIn_E[62] tile/dyn0_dataIn_E[63]
+ tile/dyn0_dataIn_E[6] tile/dyn0_dataIn_E[7] tile/dyn0_dataIn_E[8] tile/dyn0_dataIn_E[9]
+ tile/dyn0_dataIn_N[0] tile/dyn0_dataIn_N[10] tile/dyn0_dataIn_N[11] tile/dyn0_dataIn_N[12]
+ tile/dyn0_dataIn_N[13] tile/dyn0_dataIn_N[14] tile/dyn0_dataIn_N[15] tile/dyn0_dataIn_N[16]
+ tile/dyn0_dataIn_N[17] tile/dyn0_dataIn_N[18] tile/dyn0_dataIn_N[19] tile/dyn0_dataIn_N[1]
+ tile/dyn0_dataIn_N[20] tile/dyn0_dataIn_N[21] tile/dyn0_dataIn_N[22] tile/dyn0_dataIn_N[23]
+ tile/dyn0_dataIn_N[24] tile/dyn0_dataIn_N[25] tile/dyn0_dataIn_N[26] tile/dyn0_dataIn_N[27]
+ tile/dyn0_dataIn_N[28] tile/dyn0_dataIn_N[29] tile/dyn0_dataIn_N[2] tile/dyn0_dataIn_N[30]
+ tile/dyn0_dataIn_N[31] tile/dyn0_dataIn_N[32] tile/dyn0_dataIn_N[33] tile/dyn0_dataIn_N[34]
+ tile/dyn0_dataIn_N[35] tile/dyn0_dataIn_N[36] tile/dyn0_dataIn_N[37] tile/dyn0_dataIn_N[38]
+ tile/dyn0_dataIn_N[39] tile/dyn0_dataIn_N[3] tile/dyn0_dataIn_N[40] tile/dyn0_dataIn_N[41]
+ tile/dyn0_dataIn_N[42] tile/dyn0_dataIn_N[43] tile/dyn0_dataIn_N[44] tile/dyn0_dataIn_N[45]
+ tile/dyn0_dataIn_N[46] tile/dyn0_dataIn_N[47] tile/dyn0_dataIn_N[48] tile/dyn0_dataIn_N[49]
+ tile/dyn0_dataIn_N[4] tile/dyn0_dataIn_N[50] tile/dyn0_dataIn_N[51] tile/dyn0_dataIn_N[52]
+ tile/dyn0_dataIn_N[53] tile/dyn0_dataIn_N[54] tile/dyn0_dataIn_N[55] tile/dyn0_dataIn_N[56]
+ tile/dyn0_dataIn_N[57] tile/dyn0_dataIn_N[58] tile/dyn0_dataIn_N[59] tile/dyn0_dataIn_N[5]
+ tile/dyn0_dataIn_N[60] tile/dyn0_dataIn_N[61] tile/dyn0_dataIn_N[62] tile/dyn0_dataIn_N[63]
+ tile/dyn0_dataIn_N[6] tile/dyn0_dataIn_N[7] tile/dyn0_dataIn_N[8] tile/dyn0_dataIn_N[9]
+ tile/dyn0_dataIn_S[0] tile/dyn0_dataIn_S[10] tile/dyn0_dataIn_S[11] tile/dyn0_dataIn_S[12]
+ tile/dyn0_dataIn_S[13] tile/dyn0_dataIn_S[14] tile/dyn0_dataIn_S[15] tile/dyn0_dataIn_S[16]
+ tile/dyn0_dataIn_S[17] tile/dyn0_dataIn_S[18] tile/dyn0_dataIn_S[19] tile/dyn0_dataIn_S[1]
+ tile/dyn0_dataIn_S[20] tile/dyn0_dataIn_S[21] tile/dyn0_dataIn_S[22] tile/dyn0_dataIn_S[23]
+ tile/dyn0_dataIn_S[24] tile/dyn0_dataIn_S[25] tile/dyn0_dataIn_S[26] tile/dyn0_dataIn_S[27]
+ tile/dyn0_dataIn_S[28] tile/dyn0_dataIn_S[29] tile/dyn0_dataIn_S[2] tile/dyn0_dataIn_S[30]
+ tile/dyn0_dataIn_S[31] tile/dyn0_dataIn_S[32] tile/dyn0_dataIn_S[33] tile/dyn0_dataIn_S[34]
+ tile/dyn0_dataIn_S[35] tile/dyn0_dataIn_S[36] tile/dyn0_dataIn_S[37] tile/dyn0_dataIn_S[38]
+ tile/dyn0_dataIn_S[39] tile/dyn0_dataIn_S[3] tile/dyn0_dataIn_S[40] tile/dyn0_dataIn_S[41]
+ tile/dyn0_dataIn_S[42] tile/dyn0_dataIn_S[43] tile/dyn0_dataIn_S[44] tile/dyn0_dataIn_S[45]
+ tile/dyn0_dataIn_S[46] tile/dyn0_dataIn_S[47] tile/dyn0_dataIn_S[48] tile/dyn0_dataIn_S[49]
+ tile/dyn0_dataIn_S[4] tile/dyn0_dataIn_S[50] tile/dyn0_dataIn_S[51] tile/dyn0_dataIn_S[52]
+ tile/dyn0_dataIn_S[53] tile/dyn0_dataIn_S[54] tile/dyn0_dataIn_S[55] tile/dyn0_dataIn_S[56]
+ tile/dyn0_dataIn_S[57] tile/dyn0_dataIn_S[58] tile/dyn0_dataIn_S[59] tile/dyn0_dataIn_S[5]
+ tile/dyn0_dataIn_S[60] tile/dyn0_dataIn_S[61] tile/dyn0_dataIn_S[62] tile/dyn0_dataIn_S[63]
+ tile/dyn0_dataIn_S[6] tile/dyn0_dataIn_S[7] tile/dyn0_dataIn_S[8] tile/dyn0_dataIn_S[9]
+ tile/dyn0_dataIn_W[0] tile/dyn0_dataIn_W[10] tile/dyn0_dataIn_W[11] tile/dyn0_dataIn_W[12]
+ tile/dyn0_dataIn_W[13] tile/dyn0_dataIn_W[14] tile/dyn0_dataIn_W[15] tile/dyn0_dataIn_W[16]
+ tile/dyn0_dataIn_W[17] tile/dyn0_dataIn_W[18] tile/dyn0_dataIn_W[19] tile/dyn0_dataIn_W[1]
+ tile/dyn0_dataIn_W[20] tile/dyn0_dataIn_W[21] tile/dyn0_dataIn_W[22] tile/dyn0_dataIn_W[23]
+ tile/dyn0_dataIn_W[24] tile/dyn0_dataIn_W[25] tile/dyn0_dataIn_W[26] tile/dyn0_dataIn_W[27]
+ tile/dyn0_dataIn_W[28] tile/dyn0_dataIn_W[29] tile/dyn0_dataIn_W[2] tile/dyn0_dataIn_W[30]
+ tile/dyn0_dataIn_W[31] tile/dyn0_dataIn_W[32] tile/dyn0_dataIn_W[33] tile/dyn0_dataIn_W[34]
+ tile/dyn0_dataIn_W[35] tile/dyn0_dataIn_W[36] tile/dyn0_dataIn_W[37] tile/dyn0_dataIn_W[38]
+ tile/dyn0_dataIn_W[39] tile/dyn0_dataIn_W[3] tile/dyn0_dataIn_W[40] tile/dyn0_dataIn_W[41]
+ tile/dyn0_dataIn_W[42] tile/dyn0_dataIn_W[43] tile/dyn0_dataIn_W[44] tile/dyn0_dataIn_W[45]
+ tile/dyn0_dataIn_W[46] tile/dyn0_dataIn_W[47] tile/dyn0_dataIn_W[48] tile/dyn0_dataIn_W[49]
+ tile/dyn0_dataIn_W[4] tile/dyn0_dataIn_W[50] tile/dyn0_dataIn_W[51] tile/dyn0_dataIn_W[52]
+ tile/dyn0_dataIn_W[53] tile/dyn0_dataIn_W[54] tile/dyn0_dataIn_W[55] tile/dyn0_dataIn_W[56]
+ tile/dyn0_dataIn_W[57] tile/dyn0_dataIn_W[58] tile/dyn0_dataIn_W[59] tile/dyn0_dataIn_W[5]
+ tile/dyn0_dataIn_W[60] tile/dyn0_dataIn_W[61] tile/dyn0_dataIn_W[62] tile/dyn0_dataIn_W[63]
+ tile/dyn0_dataIn_W[6] tile/dyn0_dataIn_W[7] tile/dyn0_dataIn_W[8] tile/dyn0_dataIn_W[9]
+ tile/dyn0_validIn_E tile/dyn0_validIn_N tile/dyn0_validIn_S tile/dyn0_validIn_W
+ io_out[5] io_out[4] io_out[7] io_out[6] tile/dyn1_dEo[0] tile/dyn1_dEo[10] tile/dyn1_dEo[11]
+ tile/dyn1_dEo[12] tile/dyn1_dEo[13] tile/dyn1_dEo[14] tile/dyn1_dEo[15] tile/dyn1_dEo[16]
+ tile/dyn1_dEo[17] tile/dyn1_dEo[18] tile/dyn1_dEo[19] tile/dyn1_dEo[1] tile/dyn1_dEo[20]
+ tile/dyn1_dEo[21] tile/dyn1_dEo[22] tile/dyn1_dEo[23] tile/dyn1_dEo[24] tile/dyn1_dEo[25]
+ tile/dyn1_dEo[26] tile/dyn1_dEo[27] tile/dyn1_dEo[28] tile/dyn1_dEo[29] tile/dyn1_dEo[2]
+ tile/dyn1_dEo[30] tile/dyn1_dEo[31] tile/dyn1_dEo[32] tile/dyn1_dEo[33] tile/dyn1_dEo[34]
+ tile/dyn1_dEo[35] tile/dyn1_dEo[36] tile/dyn1_dEo[37] tile/dyn1_dEo[38] tile/dyn1_dEo[39]
+ tile/dyn1_dEo[3] tile/dyn1_dEo[40] tile/dyn1_dEo[41] tile/dyn1_dEo[42] tile/dyn1_dEo[43]
+ tile/dyn1_dEo[44] tile/dyn1_dEo[45] tile/dyn1_dEo[46] tile/dyn1_dEo[47] tile/dyn1_dEo[48]
+ tile/dyn1_dEo[49] tile/dyn1_dEo[4] tile/dyn1_dEo[50] tile/dyn1_dEo[51] tile/dyn1_dEo[52]
+ tile/dyn1_dEo[53] tile/dyn1_dEo[54] tile/dyn1_dEo[55] tile/dyn1_dEo[56] tile/dyn1_dEo[57]
+ tile/dyn1_dEo[58] tile/dyn1_dEo[59] tile/dyn1_dEo[5] tile/dyn1_dEo[60] tile/dyn1_dEo[61]
+ tile/dyn1_dEo[62] tile/dyn1_dEo[63] tile/dyn1_dEo[6] tile/dyn1_dEo[7] tile/dyn1_dEo[8]
+ tile/dyn1_dEo[9] io_out[9] tile/dyn1_dEo_yummy tile/dyn1_dNo[0] tile/dyn1_dNo[10]
+ tile/dyn1_dNo[11] tile/dyn1_dNo[12] tile/dyn1_dNo[13] tile/dyn1_dNo[14] tile/dyn1_dNo[15]
+ tile/dyn1_dNo[16] tile/dyn1_dNo[17] tile/dyn1_dNo[18] tile/dyn1_dNo[19] tile/dyn1_dNo[1]
+ tile/dyn1_dNo[20] tile/dyn1_dNo[21] tile/dyn1_dNo[22] tile/dyn1_dNo[23] tile/dyn1_dNo[24]
+ tile/dyn1_dNo[25] tile/dyn1_dNo[26] tile/dyn1_dNo[27] tile/dyn1_dNo[28] tile/dyn1_dNo[29]
+ tile/dyn1_dNo[2] tile/dyn1_dNo[30] tile/dyn1_dNo[31] tile/dyn1_dNo[32] tile/dyn1_dNo[33]
+ tile/dyn1_dNo[34] tile/dyn1_dNo[35] tile/dyn1_dNo[36] tile/dyn1_dNo[37] tile/dyn1_dNo[38]
+ tile/dyn1_dNo[39] tile/dyn1_dNo[3] tile/dyn1_dNo[40] tile/dyn1_dNo[41] tile/dyn1_dNo[42]
+ tile/dyn1_dNo[43] tile/dyn1_dNo[44] tile/dyn1_dNo[45] tile/dyn1_dNo[46] tile/dyn1_dNo[47]
+ tile/dyn1_dNo[48] tile/dyn1_dNo[49] tile/dyn1_dNo[4] tile/dyn1_dNo[50] tile/dyn1_dNo[51]
+ tile/dyn1_dNo[52] tile/dyn1_dNo[53] tile/dyn1_dNo[54] tile/dyn1_dNo[55] tile/dyn1_dNo[56]
+ tile/dyn1_dNo[57] tile/dyn1_dNo[58] tile/dyn1_dNo[59] tile/dyn1_dNo[5] tile/dyn1_dNo[60]
+ tile/dyn1_dNo[61] tile/dyn1_dNo[62] tile/dyn1_dNo[63] tile/dyn1_dNo[6] tile/dyn1_dNo[7]
+ tile/dyn1_dNo[8] tile/dyn1_dNo[9] io_out[8] tile/dyn1_dNo_yummy tile/dyn1_dSo[0]
+ tile/dyn1_dSo[10] tile/dyn1_dSo[11] tile/dyn1_dSo[12] tile/dyn1_dSo[13] tile/dyn1_dSo[14]
+ tile/dyn1_dSo[15] tile/dyn1_dSo[16] tile/dyn1_dSo[17] tile/dyn1_dSo[18] tile/dyn1_dSo[19]
+ tile/dyn1_dSo[1] tile/dyn1_dSo[20] tile/dyn1_dSo[21] tile/dyn1_dSo[22] tile/dyn1_dSo[23]
+ tile/dyn1_dSo[24] tile/dyn1_dSo[25] tile/dyn1_dSo[26] tile/dyn1_dSo[27] tile/dyn1_dSo[28]
+ tile/dyn1_dSo[29] tile/dyn1_dSo[2] tile/dyn1_dSo[30] tile/dyn1_dSo[31] tile/dyn1_dSo[32]
+ tile/dyn1_dSo[33] tile/dyn1_dSo[34] tile/dyn1_dSo[35] tile/dyn1_dSo[36] tile/dyn1_dSo[37]
+ tile/dyn1_dSo[38] tile/dyn1_dSo[39] tile/dyn1_dSo[3] tile/dyn1_dSo[40] tile/dyn1_dSo[41]
+ tile/dyn1_dSo[42] tile/dyn1_dSo[43] tile/dyn1_dSo[44] tile/dyn1_dSo[45] tile/dyn1_dSo[46]
+ tile/dyn1_dSo[47] tile/dyn1_dSo[48] tile/dyn1_dSo[49] tile/dyn1_dSo[4] tile/dyn1_dSo[50]
+ tile/dyn1_dSo[51] tile/dyn1_dSo[52] tile/dyn1_dSo[53] tile/dyn1_dSo[54] tile/dyn1_dSo[55]
+ tile/dyn1_dSo[56] tile/dyn1_dSo[57] tile/dyn1_dSo[58] tile/dyn1_dSo[59] tile/dyn1_dSo[5]
+ tile/dyn1_dSo[60] tile/dyn1_dSo[61] tile/dyn1_dSo[62] tile/dyn1_dSo[63] tile/dyn1_dSo[6]
+ tile/dyn1_dSo[7] tile/dyn1_dSo[8] tile/dyn1_dSo[9] io_out[11] tile/dyn1_dSo_yummy
+ tile/dyn1_dWo[0] tile/dyn1_dWo[10] tile/dyn1_dWo[11] tile/dyn1_dWo[12] tile/dyn1_dWo[13]
+ tile/dyn1_dWo[14] tile/dyn1_dWo[15] tile/dyn1_dWo[16] tile/dyn1_dWo[17] tile/dyn1_dWo[18]
+ tile/dyn1_dWo[19] tile/dyn1_dWo[1] tile/dyn1_dWo[20] tile/dyn1_dWo[21] tile/dyn1_dWo[22]
+ tile/dyn1_dWo[23] tile/dyn1_dWo[24] tile/dyn1_dWo[25] tile/dyn1_dWo[26] tile/dyn1_dWo[27]
+ tile/dyn1_dWo[28] tile/dyn1_dWo[29] tile/dyn1_dWo[2] tile/dyn1_dWo[30] tile/dyn1_dWo[31]
+ tile/dyn1_dWo[32] tile/dyn1_dWo[33] tile/dyn1_dWo[34] tile/dyn1_dWo[35] tile/dyn1_dWo[36]
+ tile/dyn1_dWo[37] tile/dyn1_dWo[38] tile/dyn1_dWo[39] tile/dyn1_dWo[3] tile/dyn1_dWo[40]
+ tile/dyn1_dWo[41] tile/dyn1_dWo[42] tile/dyn1_dWo[43] tile/dyn1_dWo[44] tile/dyn1_dWo[45]
+ tile/dyn1_dWo[46] tile/dyn1_dWo[47] tile/dyn1_dWo[48] tile/dyn1_dWo[49] tile/dyn1_dWo[4]
+ tile/dyn1_dWo[50] tile/dyn1_dWo[51] tile/dyn1_dWo[52] tile/dyn1_dWo[53] tile/dyn1_dWo[54]
+ tile/dyn1_dWo[55] tile/dyn1_dWo[56] tile/dyn1_dWo[57] tile/dyn1_dWo[58] tile/dyn1_dWo[59]
+ tile/dyn1_dWo[5] tile/dyn1_dWo[60] tile/dyn1_dWo[61] tile/dyn1_dWo[62] tile/dyn1_dWo[63]
+ tile/dyn1_dWo[6] tile/dyn1_dWo[7] tile/dyn1_dWo[8] tile/dyn1_dWo[9] io_out[10] tile/dyn1_dWo_yummy
+ tile/dyn1_dataIn_E[0] tile/dyn1_dataIn_E[10] tile/dyn1_dataIn_E[11] tile/dyn1_dataIn_E[12]
+ tile/dyn1_dataIn_E[13] tile/dyn1_dataIn_E[14] tile/dyn1_dataIn_E[15] tile/dyn1_dataIn_E[16]
+ tile/dyn1_dataIn_E[17] tile/dyn1_dataIn_E[18] tile/dyn1_dataIn_E[19] tile/dyn1_dataIn_E[1]
+ tile/dyn1_dataIn_E[20] tile/dyn1_dataIn_E[21] tile/dyn1_dataIn_E[22] tile/dyn1_dataIn_E[23]
+ tile/dyn1_dataIn_E[24] tile/dyn1_dataIn_E[25] tile/dyn1_dataIn_E[26] tile/dyn1_dataIn_E[27]
+ tile/dyn1_dataIn_E[28] tile/dyn1_dataIn_E[29] tile/dyn1_dataIn_E[2] tile/dyn1_dataIn_E[30]
+ tile/dyn1_dataIn_E[31] tile/dyn1_dataIn_E[32] tile/dyn1_dataIn_E[33] tile/dyn1_dataIn_E[34]
+ tile/dyn1_dataIn_E[35] tile/dyn1_dataIn_E[36] tile/dyn1_dataIn_E[37] tile/dyn1_dataIn_E[38]
+ tile/dyn1_dataIn_E[39] tile/dyn1_dataIn_E[3] tile/dyn1_dataIn_E[40] tile/dyn1_dataIn_E[41]
+ tile/dyn1_dataIn_E[42] tile/dyn1_dataIn_E[43] tile/dyn1_dataIn_E[44] tile/dyn1_dataIn_E[45]
+ tile/dyn1_dataIn_E[46] tile/dyn1_dataIn_E[47] tile/dyn1_dataIn_E[48] tile/dyn1_dataIn_E[49]
+ tile/dyn1_dataIn_E[4] tile/dyn1_dataIn_E[50] tile/dyn1_dataIn_E[51] tile/dyn1_dataIn_E[52]
+ tile/dyn1_dataIn_E[53] tile/dyn1_dataIn_E[54] tile/dyn1_dataIn_E[55] tile/dyn1_dataIn_E[56]
+ tile/dyn1_dataIn_E[57] tile/dyn1_dataIn_E[58] tile/dyn1_dataIn_E[59] tile/dyn1_dataIn_E[5]
+ tile/dyn1_dataIn_E[60] tile/dyn1_dataIn_E[61] tile/dyn1_dataIn_E[62] tile/dyn1_dataIn_E[63]
+ tile/dyn1_dataIn_E[6] tile/dyn1_dataIn_E[7] tile/dyn1_dataIn_E[8] tile/dyn1_dataIn_E[9]
+ tile/dyn1_dataIn_N[0] tile/dyn1_dataIn_N[10] tile/dyn1_dataIn_N[11] tile/dyn1_dataIn_N[12]
+ tile/dyn1_dataIn_N[13] tile/dyn1_dataIn_N[14] tile/dyn1_dataIn_N[15] tile/dyn1_dataIn_N[16]
+ tile/dyn1_dataIn_N[17] tile/dyn1_dataIn_N[18] tile/dyn1_dataIn_N[19] tile/dyn1_dataIn_N[1]
+ tile/dyn1_dataIn_N[20] tile/dyn1_dataIn_N[21] tile/dyn1_dataIn_N[22] tile/dyn1_dataIn_N[23]
+ tile/dyn1_dataIn_N[24] tile/dyn1_dataIn_N[25] tile/dyn1_dataIn_N[26] tile/dyn1_dataIn_N[27]
+ tile/dyn1_dataIn_N[28] tile/dyn1_dataIn_N[29] tile/dyn1_dataIn_N[2] tile/dyn1_dataIn_N[30]
+ tile/dyn1_dataIn_N[31] tile/dyn1_dataIn_N[32] tile/dyn1_dataIn_N[33] tile/dyn1_dataIn_N[34]
+ tile/dyn1_dataIn_N[35] tile/dyn1_dataIn_N[36] tile/dyn1_dataIn_N[37] tile/dyn1_dataIn_N[38]
+ tile/dyn1_dataIn_N[39] tile/dyn1_dataIn_N[3] tile/dyn1_dataIn_N[40] tile/dyn1_dataIn_N[41]
+ tile/dyn1_dataIn_N[42] tile/dyn1_dataIn_N[43] tile/dyn1_dataIn_N[44] tile/dyn1_dataIn_N[45]
+ tile/dyn1_dataIn_N[46] tile/dyn1_dataIn_N[47] tile/dyn1_dataIn_N[48] tile/dyn1_dataIn_N[49]
+ tile/dyn1_dataIn_N[4] tile/dyn1_dataIn_N[50] tile/dyn1_dataIn_N[51] tile/dyn1_dataIn_N[52]
+ tile/dyn1_dataIn_N[53] tile/dyn1_dataIn_N[54] tile/dyn1_dataIn_N[55] tile/dyn1_dataIn_N[56]
+ tile/dyn1_dataIn_N[57] tile/dyn1_dataIn_N[58] tile/dyn1_dataIn_N[59] tile/dyn1_dataIn_N[5]
+ tile/dyn1_dataIn_N[60] tile/dyn1_dataIn_N[61] tile/dyn1_dataIn_N[62] tile/dyn1_dataIn_N[63]
+ tile/dyn1_dataIn_N[6] tile/dyn1_dataIn_N[7] tile/dyn1_dataIn_N[8] tile/dyn1_dataIn_N[9]
+ tile/dyn1_dataIn_S[0] tile/dyn1_dataIn_S[10] tile/dyn1_dataIn_S[11] tile/dyn1_dataIn_S[12]
+ tile/dyn1_dataIn_S[13] tile/dyn1_dataIn_S[14] tile/dyn1_dataIn_S[15] tile/dyn1_dataIn_S[16]
+ tile/dyn1_dataIn_S[17] tile/dyn1_dataIn_S[18] tile/dyn1_dataIn_S[19] tile/dyn1_dataIn_S[1]
+ tile/dyn1_dataIn_S[20] tile/dyn1_dataIn_S[21] tile/dyn1_dataIn_S[22] tile/dyn1_dataIn_S[23]
+ tile/dyn1_dataIn_S[24] tile/dyn1_dataIn_S[25] tile/dyn1_dataIn_S[26] tile/dyn1_dataIn_S[27]
+ tile/dyn1_dataIn_S[28] tile/dyn1_dataIn_S[29] tile/dyn1_dataIn_S[2] tile/dyn1_dataIn_S[30]
+ tile/dyn1_dataIn_S[31] tile/dyn1_dataIn_S[32] tile/dyn1_dataIn_S[33] tile/dyn1_dataIn_S[34]
+ tile/dyn1_dataIn_S[35] tile/dyn1_dataIn_S[36] tile/dyn1_dataIn_S[37] tile/dyn1_dataIn_S[38]
+ tile/dyn1_dataIn_S[39] tile/dyn1_dataIn_S[3] tile/dyn1_dataIn_S[40] tile/dyn1_dataIn_S[41]
+ tile/dyn1_dataIn_S[42] tile/dyn1_dataIn_S[43] tile/dyn1_dataIn_S[44] tile/dyn1_dataIn_S[45]
+ tile/dyn1_dataIn_S[46] tile/dyn1_dataIn_S[47] tile/dyn1_dataIn_S[48] tile/dyn1_dataIn_S[49]
+ tile/dyn1_dataIn_S[4] tile/dyn1_dataIn_S[50] tile/dyn1_dataIn_S[51] tile/dyn1_dataIn_S[52]
+ tile/dyn1_dataIn_S[53] tile/dyn1_dataIn_S[54] tile/dyn1_dataIn_S[55] tile/dyn1_dataIn_S[56]
+ tile/dyn1_dataIn_S[57] tile/dyn1_dataIn_S[58] tile/dyn1_dataIn_S[59] tile/dyn1_dataIn_S[5]
+ tile/dyn1_dataIn_S[60] tile/dyn1_dataIn_S[61] tile/dyn1_dataIn_S[62] tile/dyn1_dataIn_S[63]
+ tile/dyn1_dataIn_S[6] tile/dyn1_dataIn_S[7] tile/dyn1_dataIn_S[8] tile/dyn1_dataIn_S[9]
+ tile/dyn1_dataIn_W[0] tile/dyn1_dataIn_W[10] tile/dyn1_dataIn_W[11] tile/dyn1_dataIn_W[12]
+ tile/dyn1_dataIn_W[13] tile/dyn1_dataIn_W[14] tile/dyn1_dataIn_W[15] tile/dyn1_dataIn_W[16]
+ tile/dyn1_dataIn_W[17] tile/dyn1_dataIn_W[18] tile/dyn1_dataIn_W[19] tile/dyn1_dataIn_W[1]
+ tile/dyn1_dataIn_W[20] tile/dyn1_dataIn_W[21] tile/dyn1_dataIn_W[22] tile/dyn1_dataIn_W[23]
+ tile/dyn1_dataIn_W[24] tile/dyn1_dataIn_W[25] tile/dyn1_dataIn_W[26] tile/dyn1_dataIn_W[27]
+ tile/dyn1_dataIn_W[28] tile/dyn1_dataIn_W[29] tile/dyn1_dataIn_W[2] tile/dyn1_dataIn_W[30]
+ tile/dyn1_dataIn_W[31] tile/dyn1_dataIn_W[32] tile/dyn1_dataIn_W[33] tile/dyn1_dataIn_W[34]
+ tile/dyn1_dataIn_W[35] tile/dyn1_dataIn_W[36] tile/dyn1_dataIn_W[37] tile/dyn1_dataIn_W[38]
+ tile/dyn1_dataIn_W[39] tile/dyn1_dataIn_W[3] tile/dyn1_dataIn_W[40] tile/dyn1_dataIn_W[41]
+ tile/dyn1_dataIn_W[42] tile/dyn1_dataIn_W[43] tile/dyn1_dataIn_W[44] tile/dyn1_dataIn_W[45]
+ tile/dyn1_dataIn_W[46] tile/dyn1_dataIn_W[47] tile/dyn1_dataIn_W[48] tile/dyn1_dataIn_W[49]
+ tile/dyn1_dataIn_W[4] tile/dyn1_dataIn_W[50] tile/dyn1_dataIn_W[51] tile/dyn1_dataIn_W[52]
+ tile/dyn1_dataIn_W[53] tile/dyn1_dataIn_W[54] tile/dyn1_dataIn_W[55] tile/dyn1_dataIn_W[56]
+ tile/dyn1_dataIn_W[57] tile/dyn1_dataIn_W[58] tile/dyn1_dataIn_W[59] tile/dyn1_dataIn_W[5]
+ tile/dyn1_dataIn_W[60] tile/dyn1_dataIn_W[61] tile/dyn1_dataIn_W[62] tile/dyn1_dataIn_W[63]
+ tile/dyn1_dataIn_W[6] tile/dyn1_dataIn_W[7] tile/dyn1_dataIn_W[8] tile/dyn1_dataIn_W[9]
+ tile/dyn1_validIn_E tile/dyn1_validIn_N tile/dyn1_validIn_S tile/dyn1_validIn_W
+ io_out[13] io_out[12] io_out[15] io_out[14] tile/dyn2_dEo[0] tile/dyn2_dEo[10] tile/dyn2_dEo[11]
+ tile/dyn2_dEo[12] tile/dyn2_dEo[13] tile/dyn2_dEo[14] tile/dyn2_dEo[15] tile/dyn2_dEo[16]
+ tile/dyn2_dEo[17] tile/dyn2_dEo[18] tile/dyn2_dEo[19] tile/dyn2_dEo[1] tile/dyn2_dEo[20]
+ tile/dyn2_dEo[21] tile/dyn2_dEo[22] tile/dyn2_dEo[23] tile/dyn2_dEo[24] tile/dyn2_dEo[25]
+ tile/dyn2_dEo[26] tile/dyn2_dEo[27] tile/dyn2_dEo[28] tile/dyn2_dEo[29] tile/dyn2_dEo[2]
+ tile/dyn2_dEo[30] tile/dyn2_dEo[31] tile/dyn2_dEo[32] tile/dyn2_dEo[33] tile/dyn2_dEo[34]
+ tile/dyn2_dEo[35] tile/dyn2_dEo[36] tile/dyn2_dEo[37] tile/dyn2_dEo[38] tile/dyn2_dEo[39]
+ tile/dyn2_dEo[3] tile/dyn2_dEo[40] tile/dyn2_dEo[41] tile/dyn2_dEo[42] tile/dyn2_dEo[43]
+ tile/dyn2_dEo[44] tile/dyn2_dEo[45] tile/dyn2_dEo[46] tile/dyn2_dEo[47] tile/dyn2_dEo[48]
+ tile/dyn2_dEo[49] tile/dyn2_dEo[4] tile/dyn2_dEo[50] tile/dyn2_dEo[51] tile/dyn2_dEo[52]
+ tile/dyn2_dEo[53] tile/dyn2_dEo[54] tile/dyn2_dEo[55] tile/dyn2_dEo[56] tile/dyn2_dEo[57]
+ tile/dyn2_dEo[58] tile/dyn2_dEo[59] tile/dyn2_dEo[5] tile/dyn2_dEo[60] tile/dyn2_dEo[61]
+ tile/dyn2_dEo[62] tile/dyn2_dEo[63] tile/dyn2_dEo[6] tile/dyn2_dEo[7] tile/dyn2_dEo[8]
+ tile/dyn2_dEo[9] io_out[17] tile/dyn2_dEo_yummy tile/dyn2_dNo[0] tile/dyn2_dNo[10]
+ tile/dyn2_dNo[11] tile/dyn2_dNo[12] tile/dyn2_dNo[13] tile/dyn2_dNo[14] tile/dyn2_dNo[15]
+ tile/dyn2_dNo[16] tile/dyn2_dNo[17] tile/dyn2_dNo[18] tile/dyn2_dNo[19] tile/dyn2_dNo[1]
+ tile/dyn2_dNo[20] tile/dyn2_dNo[21] tile/dyn2_dNo[22] tile/dyn2_dNo[23] tile/dyn2_dNo[24]
+ tile/dyn2_dNo[25] tile/dyn2_dNo[26] tile/dyn2_dNo[27] tile/dyn2_dNo[28] tile/dyn2_dNo[29]
+ tile/dyn2_dNo[2] tile/dyn2_dNo[30] tile/dyn2_dNo[31] tile/dyn2_dNo[32] tile/dyn2_dNo[33]
+ tile/dyn2_dNo[34] tile/dyn2_dNo[35] tile/dyn2_dNo[36] tile/dyn2_dNo[37] tile/dyn2_dNo[38]
+ tile/dyn2_dNo[39] tile/dyn2_dNo[3] tile/dyn2_dNo[40] tile/dyn2_dNo[41] tile/dyn2_dNo[42]
+ tile/dyn2_dNo[43] tile/dyn2_dNo[44] tile/dyn2_dNo[45] tile/dyn2_dNo[46] tile/dyn2_dNo[47]
+ tile/dyn2_dNo[48] tile/dyn2_dNo[49] tile/dyn2_dNo[4] tile/dyn2_dNo[50] tile/dyn2_dNo[51]
+ tile/dyn2_dNo[52] tile/dyn2_dNo[53] tile/dyn2_dNo[54] tile/dyn2_dNo[55] tile/dyn2_dNo[56]
+ tile/dyn2_dNo[57] tile/dyn2_dNo[58] tile/dyn2_dNo[59] tile/dyn2_dNo[5] tile/dyn2_dNo[60]
+ tile/dyn2_dNo[61] tile/dyn2_dNo[62] tile/dyn2_dNo[63] tile/dyn2_dNo[6] tile/dyn2_dNo[7]
+ tile/dyn2_dNo[8] tile/dyn2_dNo[9] io_out[16] tile/dyn2_dNo_yummy tile/dyn2_dSo[0]
+ tile/dyn2_dSo[10] tile/dyn2_dSo[11] tile/dyn2_dSo[12] tile/dyn2_dSo[13] tile/dyn2_dSo[14]
+ tile/dyn2_dSo[15] tile/dyn2_dSo[16] tile/dyn2_dSo[17] tile/dyn2_dSo[18] tile/dyn2_dSo[19]
+ tile/dyn2_dSo[1] tile/dyn2_dSo[20] tile/dyn2_dSo[21] tile/dyn2_dSo[22] tile/dyn2_dSo[23]
+ tile/dyn2_dSo[24] tile/dyn2_dSo[25] tile/dyn2_dSo[26] tile/dyn2_dSo[27] tile/dyn2_dSo[28]
+ tile/dyn2_dSo[29] tile/dyn2_dSo[2] tile/dyn2_dSo[30] tile/dyn2_dSo[31] tile/dyn2_dSo[32]
+ tile/dyn2_dSo[33] tile/dyn2_dSo[34] tile/dyn2_dSo[35] tile/dyn2_dSo[36] tile/dyn2_dSo[37]
+ tile/dyn2_dSo[38] tile/dyn2_dSo[39] tile/dyn2_dSo[3] tile/dyn2_dSo[40] tile/dyn2_dSo[41]
+ tile/dyn2_dSo[42] tile/dyn2_dSo[43] tile/dyn2_dSo[44] tile/dyn2_dSo[45] tile/dyn2_dSo[46]
+ tile/dyn2_dSo[47] tile/dyn2_dSo[48] tile/dyn2_dSo[49] tile/dyn2_dSo[4] tile/dyn2_dSo[50]
+ tile/dyn2_dSo[51] tile/dyn2_dSo[52] tile/dyn2_dSo[53] tile/dyn2_dSo[54] tile/dyn2_dSo[55]
+ tile/dyn2_dSo[56] tile/dyn2_dSo[57] tile/dyn2_dSo[58] tile/dyn2_dSo[59] tile/dyn2_dSo[5]
+ tile/dyn2_dSo[60] tile/dyn2_dSo[61] tile/dyn2_dSo[62] tile/dyn2_dSo[63] tile/dyn2_dSo[6]
+ tile/dyn2_dSo[7] tile/dyn2_dSo[8] tile/dyn2_dSo[9] io_out[19] tile/dyn2_dSo_yummy
+ tile/dyn2_dWo[0] tile/dyn2_dWo[10] tile/dyn2_dWo[11] tile/dyn2_dWo[12] tile/dyn2_dWo[13]
+ tile/dyn2_dWo[14] tile/dyn2_dWo[15] tile/dyn2_dWo[16] tile/dyn2_dWo[17] tile/dyn2_dWo[18]
+ tile/dyn2_dWo[19] tile/dyn2_dWo[1] tile/dyn2_dWo[20] tile/dyn2_dWo[21] tile/dyn2_dWo[22]
+ tile/dyn2_dWo[23] tile/dyn2_dWo[24] tile/dyn2_dWo[25] tile/dyn2_dWo[26] tile/dyn2_dWo[27]
+ tile/dyn2_dWo[28] tile/dyn2_dWo[29] tile/dyn2_dWo[2] tile/dyn2_dWo[30] tile/dyn2_dWo[31]
+ tile/dyn2_dWo[32] tile/dyn2_dWo[33] tile/dyn2_dWo[34] tile/dyn2_dWo[35] tile/dyn2_dWo[36]
+ tile/dyn2_dWo[37] tile/dyn2_dWo[38] tile/dyn2_dWo[39] tile/dyn2_dWo[3] tile/dyn2_dWo[40]
+ tile/dyn2_dWo[41] tile/dyn2_dWo[42] tile/dyn2_dWo[43] tile/dyn2_dWo[44] tile/dyn2_dWo[45]
+ tile/dyn2_dWo[46] tile/dyn2_dWo[47] tile/dyn2_dWo[48] tile/dyn2_dWo[49] tile/dyn2_dWo[4]
+ tile/dyn2_dWo[50] tile/dyn2_dWo[51] tile/dyn2_dWo[52] tile/dyn2_dWo[53] tile/dyn2_dWo[54]
+ tile/dyn2_dWo[55] tile/dyn2_dWo[56] tile/dyn2_dWo[57] tile/dyn2_dWo[58] tile/dyn2_dWo[59]
+ tile/dyn2_dWo[5] tile/dyn2_dWo[60] tile/dyn2_dWo[61] tile/dyn2_dWo[62] tile/dyn2_dWo[63]
+ tile/dyn2_dWo[6] tile/dyn2_dWo[7] tile/dyn2_dWo[8] tile/dyn2_dWo[9] io_out[18] tile/dyn2_dWo_yummy
+ tile/dyn2_dataIn_E[0] tile/dyn2_dataIn_E[10] tile/dyn2_dataIn_E[11] tile/dyn2_dataIn_E[12]
+ tile/dyn2_dataIn_E[13] tile/dyn2_dataIn_E[14] tile/dyn2_dataIn_E[15] tile/dyn2_dataIn_E[16]
+ tile/dyn2_dataIn_E[17] tile/dyn2_dataIn_E[18] tile/dyn2_dataIn_E[19] tile/dyn2_dataIn_E[1]
+ tile/dyn2_dataIn_E[20] tile/dyn2_dataIn_E[21] tile/dyn2_dataIn_E[22] tile/dyn2_dataIn_E[23]
+ tile/dyn2_dataIn_E[24] tile/dyn2_dataIn_E[25] tile/dyn2_dataIn_E[26] tile/dyn2_dataIn_E[27]
+ tile/dyn2_dataIn_E[28] tile/dyn2_dataIn_E[29] tile/dyn2_dataIn_E[2] tile/dyn2_dataIn_E[30]
+ tile/dyn2_dataIn_E[31] tile/dyn2_dataIn_E[32] tile/dyn2_dataIn_E[33] tile/dyn2_dataIn_E[34]
+ tile/dyn2_dataIn_E[35] tile/dyn2_dataIn_E[36] tile/dyn2_dataIn_E[37] tile/dyn2_dataIn_E[38]
+ tile/dyn2_dataIn_E[39] tile/dyn2_dataIn_E[3] tile/dyn2_dataIn_E[40] tile/dyn2_dataIn_E[41]
+ tile/dyn2_dataIn_E[42] tile/dyn2_dataIn_E[43] tile/dyn2_dataIn_E[44] tile/dyn2_dataIn_E[45]
+ tile/dyn2_dataIn_E[46] tile/dyn2_dataIn_E[47] tile/dyn2_dataIn_E[48] tile/dyn2_dataIn_E[49]
+ tile/dyn2_dataIn_E[4] tile/dyn2_dataIn_E[50] tile/dyn2_dataIn_E[51] tile/dyn2_dataIn_E[52]
+ tile/dyn2_dataIn_E[53] tile/dyn2_dataIn_E[54] tile/dyn2_dataIn_E[55] tile/dyn2_dataIn_E[56]
+ tile/dyn2_dataIn_E[57] tile/dyn2_dataIn_E[58] tile/dyn2_dataIn_E[59] tile/dyn2_dataIn_E[5]
+ tile/dyn2_dataIn_E[60] tile/dyn2_dataIn_E[61] tile/dyn2_dataIn_E[62] tile/dyn2_dataIn_E[63]
+ tile/dyn2_dataIn_E[6] tile/dyn2_dataIn_E[7] tile/dyn2_dataIn_E[8] tile/dyn2_dataIn_E[9]
+ tile/dyn2_dataIn_N[0] tile/dyn2_dataIn_N[10] tile/dyn2_dataIn_N[11] tile/dyn2_dataIn_N[12]
+ tile/dyn2_dataIn_N[13] tile/dyn2_dataIn_N[14] tile/dyn2_dataIn_N[15] tile/dyn2_dataIn_N[16]
+ tile/dyn2_dataIn_N[17] tile/dyn2_dataIn_N[18] tile/dyn2_dataIn_N[19] tile/dyn2_dataIn_N[1]
+ tile/dyn2_dataIn_N[20] tile/dyn2_dataIn_N[21] tile/dyn2_dataIn_N[22] tile/dyn2_dataIn_N[23]
+ tile/dyn2_dataIn_N[24] tile/dyn2_dataIn_N[25] tile/dyn2_dataIn_N[26] tile/dyn2_dataIn_N[27]
+ tile/dyn2_dataIn_N[28] tile/dyn2_dataIn_N[29] tile/dyn2_dataIn_N[2] tile/dyn2_dataIn_N[30]
+ tile/dyn2_dataIn_N[31] tile/dyn2_dataIn_N[32] tile/dyn2_dataIn_N[33] tile/dyn2_dataIn_N[34]
+ tile/dyn2_dataIn_N[35] tile/dyn2_dataIn_N[36] tile/dyn2_dataIn_N[37] tile/dyn2_dataIn_N[38]
+ tile/dyn2_dataIn_N[39] tile/dyn2_dataIn_N[3] tile/dyn2_dataIn_N[40] tile/dyn2_dataIn_N[41]
+ tile/dyn2_dataIn_N[42] tile/dyn2_dataIn_N[43] tile/dyn2_dataIn_N[44] tile/dyn2_dataIn_N[45]
+ tile/dyn2_dataIn_N[46] tile/dyn2_dataIn_N[47] tile/dyn2_dataIn_N[48] tile/dyn2_dataIn_N[49]
+ tile/dyn2_dataIn_N[4] tile/dyn2_dataIn_N[50] tile/dyn2_dataIn_N[51] tile/dyn2_dataIn_N[52]
+ tile/dyn2_dataIn_N[53] tile/dyn2_dataIn_N[54] tile/dyn2_dataIn_N[55] tile/dyn2_dataIn_N[56]
+ tile/dyn2_dataIn_N[57] tile/dyn2_dataIn_N[58] tile/dyn2_dataIn_N[59] tile/dyn2_dataIn_N[5]
+ tile/dyn2_dataIn_N[60] tile/dyn2_dataIn_N[61] tile/dyn2_dataIn_N[62] tile/dyn2_dataIn_N[63]
+ tile/dyn2_dataIn_N[6] tile/dyn2_dataIn_N[7] tile/dyn2_dataIn_N[8] tile/dyn2_dataIn_N[9]
+ tile/dyn2_dataIn_S[0] tile/dyn2_dataIn_S[10] tile/dyn2_dataIn_S[11] tile/dyn2_dataIn_S[12]
+ tile/dyn2_dataIn_S[13] tile/dyn2_dataIn_S[14] tile/dyn2_dataIn_S[15] tile/dyn2_dataIn_S[16]
+ tile/dyn2_dataIn_S[17] tile/dyn2_dataIn_S[18] tile/dyn2_dataIn_S[19] tile/dyn2_dataIn_S[1]
+ tile/dyn2_dataIn_S[20] tile/dyn2_dataIn_S[21] tile/dyn2_dataIn_S[22] tile/dyn2_dataIn_S[23]
+ tile/dyn2_dataIn_S[24] tile/dyn2_dataIn_S[25] tile/dyn2_dataIn_S[26] tile/dyn2_dataIn_S[27]
+ tile/dyn2_dataIn_S[28] tile/dyn2_dataIn_S[29] tile/dyn2_dataIn_S[2] tile/dyn2_dataIn_S[30]
+ tile/dyn2_dataIn_S[31] tile/dyn2_dataIn_S[32] tile/dyn2_dataIn_S[33] tile/dyn2_dataIn_S[34]
+ tile/dyn2_dataIn_S[35] tile/dyn2_dataIn_S[36] tile/dyn2_dataIn_S[37] tile/dyn2_dataIn_S[38]
+ tile/dyn2_dataIn_S[39] tile/dyn2_dataIn_S[3] tile/dyn2_dataIn_S[40] tile/dyn2_dataIn_S[41]
+ tile/dyn2_dataIn_S[42] tile/dyn2_dataIn_S[43] tile/dyn2_dataIn_S[44] tile/dyn2_dataIn_S[45]
+ tile/dyn2_dataIn_S[46] tile/dyn2_dataIn_S[47] tile/dyn2_dataIn_S[48] tile/dyn2_dataIn_S[49]
+ tile/dyn2_dataIn_S[4] tile/dyn2_dataIn_S[50] tile/dyn2_dataIn_S[51] tile/dyn2_dataIn_S[52]
+ tile/dyn2_dataIn_S[53] tile/dyn2_dataIn_S[54] tile/dyn2_dataIn_S[55] tile/dyn2_dataIn_S[56]
+ tile/dyn2_dataIn_S[57] tile/dyn2_dataIn_S[58] tile/dyn2_dataIn_S[59] tile/dyn2_dataIn_S[5]
+ tile/dyn2_dataIn_S[60] tile/dyn2_dataIn_S[61] tile/dyn2_dataIn_S[62] tile/dyn2_dataIn_S[63]
+ tile/dyn2_dataIn_S[6] tile/dyn2_dataIn_S[7] tile/dyn2_dataIn_S[8] tile/dyn2_dataIn_S[9]
+ tile/dyn2_dataIn_W[0] tile/dyn2_dataIn_W[10] tile/dyn2_dataIn_W[11] tile/dyn2_dataIn_W[12]
+ tile/dyn2_dataIn_W[13] tile/dyn2_dataIn_W[14] tile/dyn2_dataIn_W[15] tile/dyn2_dataIn_W[16]
+ tile/dyn2_dataIn_W[17] tile/dyn2_dataIn_W[18] tile/dyn2_dataIn_W[19] tile/dyn2_dataIn_W[1]
+ tile/dyn2_dataIn_W[20] tile/dyn2_dataIn_W[21] tile/dyn2_dataIn_W[22] tile/dyn2_dataIn_W[23]
+ tile/dyn2_dataIn_W[24] tile/dyn2_dataIn_W[25] tile/dyn2_dataIn_W[26] tile/dyn2_dataIn_W[27]
+ tile/dyn2_dataIn_W[28] tile/dyn2_dataIn_W[29] tile/dyn2_dataIn_W[2] tile/dyn2_dataIn_W[30]
+ tile/dyn2_dataIn_W[31] tile/dyn2_dataIn_W[32] tile/dyn2_dataIn_W[33] tile/dyn2_dataIn_W[34]
+ tile/dyn2_dataIn_W[35] tile/dyn2_dataIn_W[36] tile/dyn2_dataIn_W[37] tile/dyn2_dataIn_W[38]
+ tile/dyn2_dataIn_W[39] tile/dyn2_dataIn_W[3] tile/dyn2_dataIn_W[40] tile/dyn2_dataIn_W[41]
+ tile/dyn2_dataIn_W[42] tile/dyn2_dataIn_W[43] tile/dyn2_dataIn_W[44] tile/dyn2_dataIn_W[45]
+ tile/dyn2_dataIn_W[46] tile/dyn2_dataIn_W[47] tile/dyn2_dataIn_W[48] tile/dyn2_dataIn_W[49]
+ tile/dyn2_dataIn_W[4] tile/dyn2_dataIn_W[50] tile/dyn2_dataIn_W[51] tile/dyn2_dataIn_W[52]
+ tile/dyn2_dataIn_W[53] tile/dyn2_dataIn_W[54] tile/dyn2_dataIn_W[55] tile/dyn2_dataIn_W[56]
+ tile/dyn2_dataIn_W[57] tile/dyn2_dataIn_W[58] tile/dyn2_dataIn_W[59] tile/dyn2_dataIn_W[5]
+ tile/dyn2_dataIn_W[60] tile/dyn2_dataIn_W[61] tile/dyn2_dataIn_W[62] tile/dyn2_dataIn_W[63]
+ tile/dyn2_dataIn_W[6] tile/dyn2_dataIn_W[7] tile/dyn2_dataIn_W[8] tile/dyn2_dataIn_W[9]
+ tile/dyn2_validIn_E tile/dyn2_validIn_N tile/dyn2_validIn_S tile/dyn2_validIn_W
+ io_out[21] io_out[20] io_out[23] io_out[22] tile/flat_tileid[0] tile/flat_tileid[1]
+ tile/flat_tileid[2] tile/flat_tileid[3] tile/flat_tileid[4] tile/flat_tileid[5]
+ tile/flat_tileid[6] tile/flat_tileid[7] tile/jtag_tiles_ucb_data[0] tile/jtag_tiles_ucb_data[1]
+ tile/jtag_tiles_ucb_data[2] tile/jtag_tiles_ucb_data[3] tile/jtag_tiles_ucb_val
+ tile/l15_config_req_address_s2[10] tile/l15_config_req_address_s2[11] tile/l15_config_req_address_s2[12]
+ tile/l15_config_req_address_s2[13] tile/l15_config_req_address_s2[14] tile/l15_config_req_address_s2[15]
+ tile/l15_config_req_address_s2[8] tile/l15_config_req_address_s2[9] tile/l15_config_req_rw_s2
+ tile/l15_config_req_val_s2 tile/l15_config_write_req_data_s2[0] tile/l15_config_write_req_data_s2[10]
+ tile/l15_config_write_req_data_s2[11] tile/l15_config_write_req_data_s2[12] tile/l15_config_write_req_data_s2[13]
+ tile/l15_config_write_req_data_s2[14] tile/l15_config_write_req_data_s2[15] tile/l15_config_write_req_data_s2[16]
+ tile/l15_config_write_req_data_s2[17] tile/l15_config_write_req_data_s2[18] tile/l15_config_write_req_data_s2[19]
+ tile/l15_config_write_req_data_s2[1] tile/l15_config_write_req_data_s2[20] tile/l15_config_write_req_data_s2[21]
+ tile/l15_config_write_req_data_s2[22] tile/l15_config_write_req_data_s2[23] tile/l15_config_write_req_data_s2[24]
+ tile/l15_config_write_req_data_s2[25] tile/l15_config_write_req_data_s2[26] tile/l15_config_write_req_data_s2[27]
+ tile/l15_config_write_req_data_s2[28] tile/l15_config_write_req_data_s2[29] tile/l15_config_write_req_data_s2[2]
+ tile/l15_config_write_req_data_s2[30] tile/l15_config_write_req_data_s2[31] tile/l15_config_write_req_data_s2[32]
+ tile/l15_config_write_req_data_s2[33] tile/l15_config_write_req_data_s2[34] tile/l15_config_write_req_data_s2[35]
+ tile/l15_config_write_req_data_s2[36] tile/l15_config_write_req_data_s2[37] tile/l15_config_write_req_data_s2[38]
+ tile/l15_config_write_req_data_s2[39] tile/l15_config_write_req_data_s2[3] tile/l15_config_write_req_data_s2[40]
+ tile/l15_config_write_req_data_s2[41] tile/l15_config_write_req_data_s2[42] tile/l15_config_write_req_data_s2[43]
+ tile/l15_config_write_req_data_s2[44] tile/l15_config_write_req_data_s2[45] tile/l15_config_write_req_data_s2[46]
+ tile/l15_config_write_req_data_s2[47] tile/l15_config_write_req_data_s2[48] tile/l15_config_write_req_data_s2[49]
+ tile/l15_config_write_req_data_s2[4] tile/l15_config_write_req_data_s2[50] tile/l15_config_write_req_data_s2[51]
+ tile/l15_config_write_req_data_s2[52] tile/l15_config_write_req_data_s2[53] tile/l15_config_write_req_data_s2[54]
+ tile/l15_config_write_req_data_s2[55] tile/l15_config_write_req_data_s2[56] tile/l15_config_write_req_data_s2[57]
+ tile/l15_config_write_req_data_s2[58] tile/l15_config_write_req_data_s2[59] tile/l15_config_write_req_data_s2[5]
+ tile/l15_config_write_req_data_s2[60] tile/l15_config_write_req_data_s2[61] tile/l15_config_write_req_data_s2[62]
+ tile/l15_config_write_req_data_s2[63] tile/l15_config_write_req_data_s2[6] tile/l15_config_write_req_data_s2[7]
+ tile/l15_config_write_req_data_s2[8] tile/l15_config_write_req_data_s2[9] tile/l15_dmbr_l1missIn
+ tile/l15_dmbr_l1missTag[0] tile/l15_dmbr_l1missTag[1] tile/l15_dmbr_l1missTag[2]
+ tile/l15_dmbr_l1missTag[3] tile/l15_dmbr_l2missIn tile/l15_dmbr_l2missTag[0] tile/l15_dmbr_l2missTag[1]
+ tile/l15_dmbr_l2missTag[2] tile/l15_dmbr_l2missTag[3] tile/l15_dmbr_l2responseIn
+ tile/l15_transducer_ack tile/l15_transducer_atomic tile/l15_transducer_blockinitstore
+ tile/l15_transducer_cross_invalidate tile/l15_transducer_cross_invalidate_way[0]
+ tile/l15_transducer_cross_invalidate_way[1] tile/l15_transducer_data_0[0] tile/l15_transducer_data_0[10]
+ tile/l15_transducer_data_0[11] tile/l15_transducer_data_0[12] tile/l15_transducer_data_0[13]
+ tile/l15_transducer_data_0[14] tile/l15_transducer_data_0[15] tile/l15_transducer_data_0[16]
+ tile/l15_transducer_data_0[17] tile/l15_transducer_data_0[18] tile/l15_transducer_data_0[19]
+ tile/l15_transducer_data_0[1] tile/l15_transducer_data_0[20] tile/l15_transducer_data_0[21]
+ tile/l15_transducer_data_0[22] tile/l15_transducer_data_0[23] tile/l15_transducer_data_0[24]
+ tile/l15_transducer_data_0[25] tile/l15_transducer_data_0[26] tile/l15_transducer_data_0[27]
+ tile/l15_transducer_data_0[28] tile/l15_transducer_data_0[29] tile/l15_transducer_data_0[2]
+ tile/l15_transducer_data_0[30] tile/l15_transducer_data_0[31] tile/l15_transducer_data_0[32]
+ tile/l15_transducer_data_0[33] tile/l15_transducer_data_0[34] tile/l15_transducer_data_0[35]
+ tile/l15_transducer_data_0[36] tile/l15_transducer_data_0[37] tile/l15_transducer_data_0[38]
+ tile/l15_transducer_data_0[39] tile/l15_transducer_data_0[3] tile/l15_transducer_data_0[40]
+ tile/l15_transducer_data_0[41] tile/l15_transducer_data_0[42] tile/l15_transducer_data_0[43]
+ tile/l15_transducer_data_0[44] tile/l15_transducer_data_0[45] tile/l15_transducer_data_0[46]
+ tile/l15_transducer_data_0[47] tile/l15_transducer_data_0[48] tile/l15_transducer_data_0[49]
+ tile/l15_transducer_data_0[4] tile/l15_transducer_data_0[50] tile/l15_transducer_data_0[51]
+ tile/l15_transducer_data_0[52] tile/l15_transducer_data_0[53] tile/l15_transducer_data_0[54]
+ tile/l15_transducer_data_0[55] tile/l15_transducer_data_0[56] tile/l15_transducer_data_0[57]
+ tile/l15_transducer_data_0[58] tile/l15_transducer_data_0[59] tile/l15_transducer_data_0[5]
+ tile/l15_transducer_data_0[60] tile/l15_transducer_data_0[61] tile/l15_transducer_data_0[62]
+ tile/l15_transducer_data_0[63] tile/l15_transducer_data_0[6] tile/l15_transducer_data_0[7]
+ tile/l15_transducer_data_0[8] tile/l15_transducer_data_0[9] tile/l15_transducer_data_1[0]
+ tile/l15_transducer_data_1[10] tile/l15_transducer_data_1[11] tile/l15_transducer_data_1[12]
+ tile/l15_transducer_data_1[13] tile/l15_transducer_data_1[14] tile/l15_transducer_data_1[15]
+ tile/l15_transducer_data_1[16] tile/l15_transducer_data_1[17] tile/l15_transducer_data_1[18]
+ tile/l15_transducer_data_1[19] tile/l15_transducer_data_1[1] tile/l15_transducer_data_1[20]
+ tile/l15_transducer_data_1[21] tile/l15_transducer_data_1[22] tile/l15_transducer_data_1[23]
+ tile/l15_transducer_data_1[24] tile/l15_transducer_data_1[25] tile/l15_transducer_data_1[26]
+ tile/l15_transducer_data_1[27] tile/l15_transducer_data_1[28] tile/l15_transducer_data_1[29]
+ tile/l15_transducer_data_1[2] tile/l15_transducer_data_1[30] tile/l15_transducer_data_1[31]
+ tile/l15_transducer_data_1[32] tile/l15_transducer_data_1[33] tile/l15_transducer_data_1[34]
+ tile/l15_transducer_data_1[35] tile/l15_transducer_data_1[36] tile/l15_transducer_data_1[37]
+ tile/l15_transducer_data_1[38] tile/l15_transducer_data_1[39] tile/l15_transducer_data_1[3]
+ tile/l15_transducer_data_1[40] tile/l15_transducer_data_1[41] tile/l15_transducer_data_1[42]
+ tile/l15_transducer_data_1[43] tile/l15_transducer_data_1[44] tile/l15_transducer_data_1[45]
+ tile/l15_transducer_data_1[46] tile/l15_transducer_data_1[47] tile/l15_transducer_data_1[48]
+ tile/l15_transducer_data_1[49] tile/l15_transducer_data_1[4] tile/l15_transducer_data_1[50]
+ tile/l15_transducer_data_1[51] tile/l15_transducer_data_1[52] tile/l15_transducer_data_1[53]
+ tile/l15_transducer_data_1[54] tile/l15_transducer_data_1[55] tile/l15_transducer_data_1[56]
+ tile/l15_transducer_data_1[57] tile/l15_transducer_data_1[58] tile/l15_transducer_data_1[59]
+ tile/l15_transducer_data_1[5] tile/l15_transducer_data_1[60] tile/l15_transducer_data_1[61]
+ tile/l15_transducer_data_1[62] tile/l15_transducer_data_1[63] tile/l15_transducer_data_1[6]
+ tile/l15_transducer_data_1[7] tile/l15_transducer_data_1[8] tile/l15_transducer_data_1[9]
+ tile/l15_transducer_data_2[0] tile/l15_transducer_data_2[10] tile/l15_transducer_data_2[11]
+ tile/l15_transducer_data_2[12] tile/l15_transducer_data_2[13] tile/l15_transducer_data_2[14]
+ tile/l15_transducer_data_2[15] tile/l15_transducer_data_2[16] tile/l15_transducer_data_2[17]
+ tile/l15_transducer_data_2[18] tile/l15_transducer_data_2[19] tile/l15_transducer_data_2[1]
+ tile/l15_transducer_data_2[20] tile/l15_transducer_data_2[21] tile/l15_transducer_data_2[22]
+ tile/l15_transducer_data_2[23] tile/l15_transducer_data_2[24] tile/l15_transducer_data_2[25]
+ tile/l15_transducer_data_2[26] tile/l15_transducer_data_2[27] tile/l15_transducer_data_2[28]
+ tile/l15_transducer_data_2[29] tile/l15_transducer_data_2[2] tile/l15_transducer_data_2[30]
+ tile/l15_transducer_data_2[31] tile/l15_transducer_data_2[32] tile/l15_transducer_data_2[33]
+ tile/l15_transducer_data_2[34] tile/l15_transducer_data_2[35] tile/l15_transducer_data_2[36]
+ tile/l15_transducer_data_2[37] tile/l15_transducer_data_2[38] tile/l15_transducer_data_2[39]
+ tile/l15_transducer_data_2[3] tile/l15_transducer_data_2[40] tile/l15_transducer_data_2[41]
+ tile/l15_transducer_data_2[42] tile/l15_transducer_data_2[43] tile/l15_transducer_data_2[44]
+ tile/l15_transducer_data_2[45] tile/l15_transducer_data_2[46] tile/l15_transducer_data_2[47]
+ tile/l15_transducer_data_2[48] tile/l15_transducer_data_2[49] tile/l15_transducer_data_2[4]
+ tile/l15_transducer_data_2[50] tile/l15_transducer_data_2[51] tile/l15_transducer_data_2[52]
+ tile/l15_transducer_data_2[53] tile/l15_transducer_data_2[54] tile/l15_transducer_data_2[55]
+ tile/l15_transducer_data_2[56] tile/l15_transducer_data_2[57] tile/l15_transducer_data_2[58]
+ tile/l15_transducer_data_2[59] tile/l15_transducer_data_2[5] tile/l15_transducer_data_2[60]
+ tile/l15_transducer_data_2[61] tile/l15_transducer_data_2[62] tile/l15_transducer_data_2[63]
+ tile/l15_transducer_data_2[6] tile/l15_transducer_data_2[7] tile/l15_transducer_data_2[8]
+ tile/l15_transducer_data_2[9] tile/l15_transducer_data_3[0] tile/l15_transducer_data_3[10]
+ tile/l15_transducer_data_3[11] tile/l15_transducer_data_3[12] tile/l15_transducer_data_3[13]
+ tile/l15_transducer_data_3[14] tile/l15_transducer_data_3[15] tile/l15_transducer_data_3[16]
+ tile/l15_transducer_data_3[17] tile/l15_transducer_data_3[18] tile/l15_transducer_data_3[19]
+ tile/l15_transducer_data_3[1] tile/l15_transducer_data_3[20] tile/l15_transducer_data_3[21]
+ tile/l15_transducer_data_3[22] tile/l15_transducer_data_3[23] tile/l15_transducer_data_3[24]
+ tile/l15_transducer_data_3[25] tile/l15_transducer_data_3[26] tile/l15_transducer_data_3[27]
+ tile/l15_transducer_data_3[28] tile/l15_transducer_data_3[29] tile/l15_transducer_data_3[2]
+ tile/l15_transducer_data_3[30] tile/l15_transducer_data_3[31] tile/l15_transducer_data_3[32]
+ tile/l15_transducer_data_3[33] tile/l15_transducer_data_3[34] tile/l15_transducer_data_3[35]
+ tile/l15_transducer_data_3[36] tile/l15_transducer_data_3[37] tile/l15_transducer_data_3[38]
+ tile/l15_transducer_data_3[39] tile/l15_transducer_data_3[3] tile/l15_transducer_data_3[40]
+ tile/l15_transducer_data_3[41] tile/l15_transducer_data_3[42] tile/l15_transducer_data_3[43]
+ tile/l15_transducer_data_3[44] tile/l15_transducer_data_3[45] tile/l15_transducer_data_3[46]
+ tile/l15_transducer_data_3[47] tile/l15_transducer_data_3[48] tile/l15_transducer_data_3[49]
+ tile/l15_transducer_data_3[4] tile/l15_transducer_data_3[50] tile/l15_transducer_data_3[51]
+ tile/l15_transducer_data_3[52] tile/l15_transducer_data_3[53] tile/l15_transducer_data_3[54]
+ tile/l15_transducer_data_3[55] tile/l15_transducer_data_3[56] tile/l15_transducer_data_3[57]
+ tile/l15_transducer_data_3[58] tile/l15_transducer_data_3[59] tile/l15_transducer_data_3[5]
+ tile/l15_transducer_data_3[60] tile/l15_transducer_data_3[61] tile/l15_transducer_data_3[62]
+ tile/l15_transducer_data_3[63] tile/l15_transducer_data_3[6] tile/l15_transducer_data_3[7]
+ tile/l15_transducer_data_3[8] tile/l15_transducer_data_3[9] tile/l15_transducer_error[0]
+ tile/l15_transducer_error[1] tile/l15_transducer_f4b tile/l15_transducer_header_ack
+ tile/l15_transducer_inval_address_15_4[10] tile/l15_transducer_inval_address_15_4[11]
+ tile/l15_transducer_inval_address_15_4[12] tile/l15_transducer_inval_address_15_4[13]
+ tile/l15_transducer_inval_address_15_4[14] tile/l15_transducer_inval_address_15_4[15]
+ tile/l15_transducer_inval_address_15_4[4] tile/l15_transducer_inval_address_15_4[5]
+ tile/l15_transducer_inval_address_15_4[6] tile/l15_transducer_inval_address_15_4[7]
+ tile/l15_transducer_inval_address_15_4[8] tile/l15_transducer_inval_address_15_4[9]
+ tile/l15_transducer_inval_dcache_all_way tile/l15_transducer_inval_dcache_inval
+ tile/l15_transducer_inval_icache_all_way tile/l15_transducer_inval_icache_inval
+ tile/l15_transducer_inval_way[0] tile/l15_transducer_inval_way[1] tile/l15_transducer_l2miss
+ tile/l15_transducer_noncacheable tile/l15_transducer_prefetch tile/l15_transducer_returntype[0]
+ tile/l15_transducer_returntype[1] tile/l15_transducer_returntype[2] tile/l15_transducer_returntype[3]
+ tile/l15_transducer_threadid tile/l15_transducer_val tile/l2_rtap_data[0] tile/l2_rtap_data[1]
+ tile/l2_rtap_data[2] tile/l2_rtap_data[3] tile/noc1_out_data[0] tile/noc1_out_data[10]
+ tile/noc1_out_data[11] tile/noc1_out_data[12] tile/noc1_out_data[13] tile/noc1_out_data[14]
+ tile/noc1_out_data[15] tile/noc1_out_data[16] tile/noc1_out_data[17] tile/noc1_out_data[18]
+ tile/noc1_out_data[19] tile/noc1_out_data[1] tile/noc1_out_data[20] tile/noc1_out_data[21]
+ tile/noc1_out_data[22] tile/noc1_out_data[23] tile/noc1_out_data[24] tile/noc1_out_data[25]
+ tile/noc1_out_data[26] tile/noc1_out_data[27] tile/noc1_out_data[28] tile/noc1_out_data[29]
+ tile/noc1_out_data[2] tile/noc1_out_data[30] tile/noc1_out_data[31] tile/noc1_out_data[32]
+ tile/noc1_out_data[33] tile/noc1_out_data[34] tile/noc1_out_data[35] tile/noc1_out_data[36]
+ tile/noc1_out_data[37] tile/noc1_out_data[38] tile/noc1_out_data[39] tile/noc1_out_data[3]
+ tile/noc1_out_data[40] tile/noc1_out_data[41] tile/noc1_out_data[42] tile/noc1_out_data[43]
+ tile/noc1_out_data[44] tile/noc1_out_data[45] tile/noc1_out_data[46] tile/noc1_out_data[47]
+ tile/noc1_out_data[48] tile/noc1_out_data[49] tile/noc1_out_data[4] tile/noc1_out_data[50]
+ tile/noc1_out_data[51] tile/noc1_out_data[52] tile/noc1_out_data[53] tile/noc1_out_data[54]
+ tile/noc1_out_data[55] tile/noc1_out_data[56] tile/noc1_out_data[57] tile/noc1_out_data[58]
+ tile/noc1_out_data[59] tile/noc1_out_data[5] tile/noc1_out_data[60] tile/noc1_out_data[61]
+ tile/noc1_out_data[62] tile/noc1_out_data[63] tile/noc1_out_data[6] tile/noc1_out_data[7]
+ tile/noc1_out_data[8] tile/noc1_out_data[9] tile/noc1_out_rdy tile/noc1_out_val
+ tile/noc2_in_data[0] tile/noc2_in_data[10] tile/noc2_in_data[11] tile/noc2_in_data[12]
+ tile/noc2_in_data[13] tile/noc2_in_data[14] tile/noc2_in_data[15] tile/noc2_in_data[16]
+ tile/noc2_in_data[17] tile/noc2_in_data[18] tile/noc2_in_data[19] tile/noc2_in_data[1]
+ tile/noc2_in_data[20] tile/noc2_in_data[21] tile/noc2_in_data[22] tile/noc2_in_data[23]
+ tile/noc2_in_data[24] tile/noc2_in_data[25] tile/noc2_in_data[26] tile/noc2_in_data[27]
+ tile/noc2_in_data[28] tile/noc2_in_data[29] tile/noc2_in_data[2] tile/noc2_in_data[30]
+ tile/noc2_in_data[31] tile/noc2_in_data[32] tile/noc2_in_data[33] tile/noc2_in_data[34]
+ tile/noc2_in_data[35] tile/noc2_in_data[36] tile/noc2_in_data[37] tile/noc2_in_data[38]
+ tile/noc2_in_data[39] tile/noc2_in_data[3] tile/noc2_in_data[40] tile/noc2_in_data[41]
+ tile/noc2_in_data[42] tile/noc2_in_data[43] tile/noc2_in_data[44] tile/noc2_in_data[45]
+ tile/noc2_in_data[46] tile/noc2_in_data[47] tile/noc2_in_data[48] tile/noc2_in_data[49]
+ tile/noc2_in_data[4] tile/noc2_in_data[50] tile/noc2_in_data[51] tile/noc2_in_data[52]
+ tile/noc2_in_data[53] tile/noc2_in_data[54] tile/noc2_in_data[55] tile/noc2_in_data[56]
+ tile/noc2_in_data[57] tile/noc2_in_data[58] tile/noc2_in_data[59] tile/noc2_in_data[5]
+ tile/noc2_in_data[60] tile/noc2_in_data[61] tile/noc2_in_data[62] tile/noc2_in_data[63]
+ tile/noc2_in_data[6] tile/noc2_in_data[7] tile/noc2_in_data[8] tile/noc2_in_data[9]
+ tile/noc2_in_rdy tile/noc2_in_val tile/noc3_out_data[0] tile/noc3_out_data[10] tile/noc3_out_data[11]
+ tile/noc3_out_data[12] tile/noc3_out_data[13] tile/noc3_out_data[14] tile/noc3_out_data[15]
+ tile/noc3_out_data[16] tile/noc3_out_data[17] tile/noc3_out_data[18] tile/noc3_out_data[19]
+ tile/noc3_out_data[1] tile/noc3_out_data[20] tile/noc3_out_data[21] tile/noc3_out_data[22]
+ tile/noc3_out_data[23] tile/noc3_out_data[24] tile/noc3_out_data[25] tile/noc3_out_data[26]
+ tile/noc3_out_data[27] tile/noc3_out_data[28] tile/noc3_out_data[29] tile/noc3_out_data[2]
+ tile/noc3_out_data[30] tile/noc3_out_data[31] tile/noc3_out_data[32] tile/noc3_out_data[33]
+ tile/noc3_out_data[34] tile/noc3_out_data[35] tile/noc3_out_data[36] tile/noc3_out_data[37]
+ tile/noc3_out_data[38] tile/noc3_out_data[39] tile/noc3_out_data[3] tile/noc3_out_data[40]
+ tile/noc3_out_data[41] tile/noc3_out_data[42] tile/noc3_out_data[43] tile/noc3_out_data[44]
+ tile/noc3_out_data[45] tile/noc3_out_data[46] tile/noc3_out_data[47] tile/noc3_out_data[48]
+ tile/noc3_out_data[49] tile/noc3_out_data[4] tile/noc3_out_data[50] tile/noc3_out_data[51]
+ tile/noc3_out_data[52] tile/noc3_out_data[53] tile/noc3_out_data[54] tile/noc3_out_data[55]
+ tile/noc3_out_data[56] tile/noc3_out_data[57] tile/noc3_out_data[58] tile/noc3_out_data[59]
+ tile/noc3_out_data[5] tile/noc3_out_data[60] tile/noc3_out_data[61] tile/noc3_out_data[62]
+ tile/noc3_out_data[63] tile/noc3_out_data[6] tile/noc3_out_data[7] tile/noc3_out_data[8]
+ tile/noc3_out_data[9] tile/noc3_out_rdy tile/noc3_out_val tile/processor_router_data_noc2[0]
+ tile/processor_router_data_noc2[10] tile/processor_router_data_noc2[11] tile/processor_router_data_noc2[12]
+ tile/processor_router_data_noc2[13] tile/processor_router_data_noc2[14] tile/processor_router_data_noc2[15]
+ tile/processor_router_data_noc2[16] tile/processor_router_data_noc2[17] tile/processor_router_data_noc2[18]
+ tile/processor_router_data_noc2[19] tile/processor_router_data_noc2[1] tile/processor_router_data_noc2[20]
+ tile/processor_router_data_noc2[21] tile/processor_router_data_noc2[22] tile/processor_router_data_noc2[23]
+ tile/processor_router_data_noc2[24] tile/processor_router_data_noc2[25] tile/processor_router_data_noc2[26]
+ tile/processor_router_data_noc2[27] tile/processor_router_data_noc2[28] tile/processor_router_data_noc2[29]
+ tile/processor_router_data_noc2[2] tile/processor_router_data_noc2[30] tile/processor_router_data_noc2[31]
+ tile/processor_router_data_noc2[32] tile/processor_router_data_noc2[33] tile/processor_router_data_noc2[34]
+ tile/processor_router_data_noc2[35] tile/processor_router_data_noc2[36] tile/processor_router_data_noc2[37]
+ tile/processor_router_data_noc2[38] tile/processor_router_data_noc2[39] tile/processor_router_data_noc2[3]
+ tile/processor_router_data_noc2[40] tile/processor_router_data_noc2[41] tile/processor_router_data_noc2[42]
+ tile/processor_router_data_noc2[43] tile/processor_router_data_noc2[44] tile/processor_router_data_noc2[45]
+ tile/processor_router_data_noc2[46] tile/processor_router_data_noc2[47] tile/processor_router_data_noc2[48]
+ tile/processor_router_data_noc2[49] tile/processor_router_data_noc2[4] tile/processor_router_data_noc2[50]
+ tile/processor_router_data_noc2[51] tile/processor_router_data_noc2[52] tile/processor_router_data_noc2[53]
+ tile/processor_router_data_noc2[54] tile/processor_router_data_noc2[55] tile/processor_router_data_noc2[56]
+ tile/processor_router_data_noc2[57] tile/processor_router_data_noc2[58] tile/processor_router_data_noc2[59]
+ tile/processor_router_data_noc2[5] tile/processor_router_data_noc2[60] tile/processor_router_data_noc2[61]
+ tile/processor_router_data_noc2[62] tile/processor_router_data_noc2[63] tile/processor_router_data_noc2[6]
+ tile/processor_router_data_noc2[7] tile/processor_router_data_noc2[8] tile/processor_router_data_noc2[9]
+ tile/processor_router_ready_noc1 tile/processor_router_ready_noc3 tile/processor_router_valid_noc2
+ tile/router_processor_ready_noc2 wb_rst_i tile/rtap_srams_bist_command[0] tile/rtap_srams_bist_command[1]
+ tile/rtap_srams_bist_command[2] tile/rtap_srams_bist_command[3] tile/rtap_srams_bist_data[0]
+ tile/rtap_srams_bist_data[1] tile/rtap_srams_bist_data[2] tile/rtap_srams_bist_data[3]
+ tile/srams_rtap_data[0] tile/srams_rtap_data[1] tile/srams_rtap_data[2] tile/srams_rtap_data[3]
+ tile/tile_jtag_ucb_data[0] tile/tile_jtag_ucb_data[1] tile/tile_jtag_ucb_data[2]
+ tile/tile_jtag_ucb_data[3] tile/tile_jtag_ucb_val tile/transducer_l15_address[0]
+ tile/transducer_l15_address[10] tile/transducer_l15_address[11] tile/transducer_l15_address[12]
+ tile/transducer_l15_address[13] tile/transducer_l15_address[14] tile/transducer_l15_address[15]
+ tile/transducer_l15_address[16] tile/transducer_l15_address[17] tile/transducer_l15_address[18]
+ tile/transducer_l15_address[19] tile/transducer_l15_address[1] tile/transducer_l15_address[20]
+ tile/transducer_l15_address[21] tile/transducer_l15_address[22] tile/transducer_l15_address[23]
+ tile/transducer_l15_address[24] tile/transducer_l15_address[25] tile/transducer_l15_address[26]
+ tile/transducer_l15_address[27] tile/transducer_l15_address[28] tile/transducer_l15_address[29]
+ tile/transducer_l15_address[2] tile/transducer_l15_address[30] tile/transducer_l15_address[31]
+ tile/transducer_l15_address[32] tile/transducer_l15_address[33] tile/transducer_l15_address[34]
+ tile/transducer_l15_address[35] tile/transducer_l15_address[36] tile/transducer_l15_address[37]
+ tile/transducer_l15_address[38] tile/transducer_l15_address[39] tile/transducer_l15_address[3]
+ tile/transducer_l15_address[4] tile/transducer_l15_address[5] tile/transducer_l15_address[6]
+ tile/transducer_l15_address[7] tile/transducer_l15_address[8] tile/transducer_l15_address[9]
+ tile/transducer_l15_amo_op[0] tile/transducer_l15_amo_op[1] tile/transducer_l15_amo_op[2]
+ tile/transducer_l15_amo_op[3] tile/transducer_l15_blockinitstore tile/transducer_l15_blockstore
+ tile/transducer_l15_csm_data[0] tile/transducer_l15_csm_data[10] tile/transducer_l15_csm_data[11]
+ tile/transducer_l15_csm_data[12] tile/transducer_l15_csm_data[13] tile/transducer_l15_csm_data[14]
+ tile/transducer_l15_csm_data[15] tile/transducer_l15_csm_data[16] tile/transducer_l15_csm_data[17]
+ tile/transducer_l15_csm_data[18] tile/transducer_l15_csm_data[19] tile/transducer_l15_csm_data[1]
+ tile/transducer_l15_csm_data[20] tile/transducer_l15_csm_data[21] tile/transducer_l15_csm_data[22]
+ tile/transducer_l15_csm_data[23] tile/transducer_l15_csm_data[24] tile/transducer_l15_csm_data[25]
+ tile/transducer_l15_csm_data[26] tile/transducer_l15_csm_data[27] tile/transducer_l15_csm_data[28]
+ tile/transducer_l15_csm_data[29] tile/transducer_l15_csm_data[2] tile/transducer_l15_csm_data[30]
+ tile/transducer_l15_csm_data[31] tile/transducer_l15_csm_data[32] tile/transducer_l15_csm_data[3]
+ tile/transducer_l15_csm_data[4] tile/transducer_l15_csm_data[5] tile/transducer_l15_csm_data[6]
+ tile/transducer_l15_csm_data[7] tile/transducer_l15_csm_data[8] tile/transducer_l15_csm_data[9]
+ tile/transducer_l15_data[0] tile/transducer_l15_data[10] tile/transducer_l15_data[11]
+ tile/transducer_l15_data[12] tile/transducer_l15_data[13] tile/transducer_l15_data[14]
+ tile/transducer_l15_data[15] tile/transducer_l15_data[16] tile/transducer_l15_data[17]
+ tile/transducer_l15_data[18] tile/transducer_l15_data[19] tile/transducer_l15_data[1]
+ tile/transducer_l15_data[20] tile/transducer_l15_data[21] tile/transducer_l15_data[22]
+ tile/transducer_l15_data[23] tile/transducer_l15_data[24] tile/transducer_l15_data[25]
+ tile/transducer_l15_data[26] tile/transducer_l15_data[27] tile/transducer_l15_data[28]
+ tile/transducer_l15_data[29] tile/transducer_l15_data[2] tile/transducer_l15_data[30]
+ tile/transducer_l15_data[31] tile/transducer_l15_data[32] tile/transducer_l15_data[33]
+ tile/transducer_l15_data[34] tile/transducer_l15_data[35] tile/transducer_l15_data[36]
+ tile/transducer_l15_data[37] tile/transducer_l15_data[38] tile/transducer_l15_data[39]
+ tile/transducer_l15_data[3] tile/transducer_l15_data[40] tile/transducer_l15_data[41]
+ tile/transducer_l15_data[42] tile/transducer_l15_data[43] tile/transducer_l15_data[44]
+ tile/transducer_l15_data[45] tile/transducer_l15_data[46] tile/transducer_l15_data[47]
+ tile/transducer_l15_data[48] tile/transducer_l15_data[49] tile/transducer_l15_data[4]
+ tile/transducer_l15_data[50] tile/transducer_l15_data[51] tile/transducer_l15_data[52]
+ tile/transducer_l15_data[53] tile/transducer_l15_data[54] tile/transducer_l15_data[55]
+ tile/transducer_l15_data[56] tile/transducer_l15_data[57] tile/transducer_l15_data[58]
+ tile/transducer_l15_data[59] tile/transducer_l15_data[5] tile/transducer_l15_data[60]
+ tile/transducer_l15_data[61] tile/transducer_l15_data[62] tile/transducer_l15_data[63]
+ tile/transducer_l15_data[6] tile/transducer_l15_data[7] tile/transducer_l15_data[8]
+ tile/transducer_l15_data[9] tile/transducer_l15_data_next_entry[0] tile/transducer_l15_data_next_entry[10]
+ tile/transducer_l15_data_next_entry[11] tile/transducer_l15_data_next_entry[12]
+ tile/transducer_l15_data_next_entry[13] tile/transducer_l15_data_next_entry[14]
+ tile/transducer_l15_data_next_entry[15] tile/transducer_l15_data_next_entry[16]
+ tile/transducer_l15_data_next_entry[17] tile/transducer_l15_data_next_entry[18]
+ tile/transducer_l15_data_next_entry[19] tile/transducer_l15_data_next_entry[1] tile/transducer_l15_data_next_entry[20]
+ tile/transducer_l15_data_next_entry[21] tile/transducer_l15_data_next_entry[22]
+ tile/transducer_l15_data_next_entry[23] tile/transducer_l15_data_next_entry[24]
+ tile/transducer_l15_data_next_entry[25] tile/transducer_l15_data_next_entry[26]
+ tile/transducer_l15_data_next_entry[27] tile/transducer_l15_data_next_entry[28]
+ tile/transducer_l15_data_next_entry[29] tile/transducer_l15_data_next_entry[2] tile/transducer_l15_data_next_entry[30]
+ tile/transducer_l15_data_next_entry[31] tile/transducer_l15_data_next_entry[32]
+ tile/transducer_l15_data_next_entry[33] tile/transducer_l15_data_next_entry[34]
+ tile/transducer_l15_data_next_entry[35] tile/transducer_l15_data_next_entry[36]
+ tile/transducer_l15_data_next_entry[37] tile/transducer_l15_data_next_entry[38]
+ tile/transducer_l15_data_next_entry[39] tile/transducer_l15_data_next_entry[3] tile/transducer_l15_data_next_entry[40]
+ tile/transducer_l15_data_next_entry[41] tile/transducer_l15_data_next_entry[42]
+ tile/transducer_l15_data_next_entry[43] tile/transducer_l15_data_next_entry[44]
+ tile/transducer_l15_data_next_entry[45] tile/transducer_l15_data_next_entry[46]
+ tile/transducer_l15_data_next_entry[47] tile/transducer_l15_data_next_entry[48]
+ tile/transducer_l15_data_next_entry[49] tile/transducer_l15_data_next_entry[4] tile/transducer_l15_data_next_entry[50]
+ tile/transducer_l15_data_next_entry[51] tile/transducer_l15_data_next_entry[52]
+ tile/transducer_l15_data_next_entry[53] tile/transducer_l15_data_next_entry[54]
+ tile/transducer_l15_data_next_entry[55] tile/transducer_l15_data_next_entry[56]
+ tile/transducer_l15_data_next_entry[57] tile/transducer_l15_data_next_entry[58]
+ tile/transducer_l15_data_next_entry[59] tile/transducer_l15_data_next_entry[5] tile/transducer_l15_data_next_entry[60]
+ tile/transducer_l15_data_next_entry[61] tile/transducer_l15_data_next_entry[62]
+ tile/transducer_l15_data_next_entry[63] tile/transducer_l15_data_next_entry[6] tile/transducer_l15_data_next_entry[7]
+ tile/transducer_l15_data_next_entry[8] tile/transducer_l15_data_next_entry[9] tile/transducer_l15_invalidate_cacheline
+ tile/transducer_l15_l1rplway[0] tile/transducer_l15_l1rplway[1] tile/transducer_l15_nc
+ tile/transducer_l15_prefetch tile/transducer_l15_req_ack tile/transducer_l15_rqtype[0]
+ tile/transducer_l15_rqtype[1] tile/transducer_l15_rqtype[2] tile/transducer_l15_rqtype[3]
+ tile/transducer_l15_rqtype[4] tile/transducer_l15_size[0] tile/transducer_l15_size[1]
+ tile/transducer_l15_size[2] tile/transducer_l15_threadid tile/transducer_l15_val
+ tile/vccd1 tile/vssd1 tile
.ends

